##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Fri Jun  3 01:22:46 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO soc_now_caravel_top
  CLASS BLOCK ;
  SIZE 1420.020000 BY 1419.840000 ;
  FOREIGN soc_now_caravel_top 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 482.160000 1419.040000 482.460000 1419.840000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 490.900000 1419.040000 491.200000 1419.840000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1410.440000 1419.040000 1410.740000 1419.840000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.500000 1419.040000 794.800000 1419.840000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.640000 1419.040000 1419.940000 1419.840000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1401.700000 1419.040000 1402.000000 1419.840000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1392.500000 1419.040000 1392.800000 1419.840000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1383.760000 1419.040000 1384.060000 1419.840000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1374.560000 1419.040000 1374.860000 1419.840000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1080.160000 1419.040000 1080.460000 1419.840000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1071.420000 1419.040000 1071.720000 1419.840000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1062.220000 1419.040000 1062.520000 1419.840000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1053.480000 1419.040000 1053.780000 1419.840000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1044.280000 1419.040000 1044.580000 1419.840000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1035.540000 1419.040000 1035.840000 1419.840000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1026.800000 1419.040000 1027.100000 1419.840000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1017.600000 1419.040000 1017.900000 1419.840000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1008.860000 1419.040000 1009.160000 1419.840000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 999.660000 1419.040000 999.960000 1419.840000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 990.920000 1419.040000 991.220000 1419.840000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 981.720000 1419.040000 982.020000 1419.840000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 972.980000 1419.040000 973.280000 1419.840000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 964.240000 1419.040000 964.540000 1419.840000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 955.040000 1419.040000 955.340000 1419.840000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 946.300000 1419.040000 946.600000 1419.840000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 937.100000 1419.040000 937.400000 1419.840000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.360000 1419.040000 928.660000 1419.840000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 919.620000 1419.040000 919.920000 1419.840000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 910.420000 1419.040000 910.720000 1419.840000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 901.680000 1419.040000 901.980000 1419.840000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 892.480000 1419.040000 892.780000 1419.840000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 883.740000 1419.040000 884.040000 1419.840000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 875.000000 1419.040000 875.300000 1419.840000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 865.800000 1419.040000 866.100000 1419.840000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 857.060000 1419.040000 857.360000 1419.840000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 847.860000 1419.040000 848.160000 1419.840000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 839.120000 1419.040000 839.420000 1419.840000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 830.380000 1419.040000 830.680000 1419.840000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.180000 1419.040000 821.480000 1419.840000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 812.440000 1419.040000 812.740000 1419.840000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 803.240000 1419.040000 803.540000 1419.840000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 785.300000 1419.040000 785.600000 1419.840000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 776.560000 1419.040000 776.860000 1419.840000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 767.820000 1419.040000 768.120000 1419.840000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 758.620000 1419.040000 758.920000 1419.840000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 749.880000 1419.040000 750.180000 1419.840000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 740.680000 1419.040000 740.980000 1419.840000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 731.940000 1419.040000 732.240000 1419.840000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 723.200000 1419.040000 723.500000 1419.840000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 714.000000 1419.040000 714.300000 1419.840000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 705.260000 1419.040000 705.560000 1419.840000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.060000 1419.040000 696.360000 1419.840000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 687.320000 1419.040000 687.620000 1419.840000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 678.580000 1419.040000 678.880000 1419.840000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.380000 1419.040000 669.680000 1419.840000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 660.640000 1419.040000 660.940000 1419.840000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 651.440000 1419.040000 651.740000 1419.840000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 642.700000 1419.040000 643.000000 1419.840000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 633.960000 1419.040000 634.260000 1419.840000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 624.760000 1419.040000 625.060000 1419.840000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 616.020000 1419.040000 616.320000 1419.840000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 606.820000 1419.040000 607.120000 1419.840000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 598.080000 1419.040000 598.380000 1419.840000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 588.880000 1419.040000 589.180000 1419.840000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 580.140000 1419.040000 580.440000 1419.840000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 571.400000 1419.040000 571.700000 1419.840000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 562.200000 1419.040000 562.500000 1419.840000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 553.460000 1419.040000 553.760000 1419.840000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 544.260000 1419.040000 544.560000 1419.840000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 535.520000 1419.040000 535.820000 1419.840000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 526.780000 1419.040000 527.080000 1419.840000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 517.580000 1419.040000 517.880000 1419.840000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 508.840000 1419.040000 509.140000 1419.840000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 499.640000 1419.040000 499.940000 1419.840000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1365.820000 1419.040000 1366.120000 1419.840000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.080000 1419.040000 1357.380000 1419.840000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1347.880000 1419.040000 1348.180000 1419.840000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1339.140000 1419.040000 1339.440000 1419.840000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1329.940000 1419.040000 1330.240000 1419.840000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1321.200000 1419.040000 1321.500000 1419.840000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1312.460000 1419.040000 1312.760000 1419.840000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1303.260000 1419.040000 1303.560000 1419.840000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1294.520000 1419.040000 1294.820000 1419.840000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1285.320000 1419.040000 1285.620000 1419.840000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1276.580000 1419.040000 1276.880000 1419.840000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1267.840000 1419.040000 1268.140000 1419.840000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1258.640000 1419.040000 1258.940000 1419.840000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1249.900000 1419.040000 1250.200000 1419.840000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1240.700000 1419.040000 1241.000000 1419.840000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1231.960000 1419.040000 1232.260000 1419.840000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1223.220000 1419.040000 1223.520000 1419.840000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1214.020000 1419.040000 1214.320000 1419.840000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1205.280000 1419.040000 1205.580000 1419.840000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.080000 1419.040000 1196.380000 1419.840000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1187.340000 1419.040000 1187.640000 1419.840000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1178.140000 1419.040000 1178.440000 1419.840000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1169.400000 1419.040000 1169.700000 1419.840000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1160.660000 1419.040000 1160.960000 1419.840000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1151.460000 1419.040000 1151.760000 1419.840000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1142.720000 1419.040000 1143.020000 1419.840000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1133.520000 1419.040000 1133.820000 1419.840000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1124.780000 1419.040000 1125.080000 1419.840000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1116.040000 1419.040000 1116.340000 1419.840000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1106.840000 1419.040000 1107.140000 1419.840000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1098.100000 1419.040000 1098.400000 1419.840000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1088.900000 1419.040000 1089.200000 1419.840000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 472.960000 1419.040000 473.260000 1419.840000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 464.220000 1419.040000 464.520000 1419.840000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 455.020000 1419.040000 455.320000 1419.840000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.280000 1419.040000 446.580000 1419.840000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 437.540000 1419.040000 437.840000 1419.840000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.340000 1419.040000 428.640000 1419.840000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 419.600000 1419.040000 419.900000 1419.840000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 410.400000 1419.040000 410.700000 1419.840000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 401.660000 1419.040000 401.960000 1419.840000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 392.460000 1419.040000 392.760000 1419.840000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.720000 1419.040000 384.020000 1419.840000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 374.980000 1419.040000 375.280000 1419.840000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 365.780000 1419.040000 366.080000 1419.840000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 357.040000 1419.040000 357.340000 1419.840000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 347.840000 1419.040000 348.140000 1419.840000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 339.100000 1419.040000 339.400000 1419.840000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 330.360000 1419.040000 330.660000 1419.840000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 321.160000 1419.040000 321.460000 1419.840000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 312.420000 1419.040000 312.720000 1419.840000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 303.220000 1419.040000 303.520000 1419.840000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 294.480000 1419.040000 294.780000 1419.840000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 285.740000 1419.040000 286.040000 1419.840000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 276.540000 1419.040000 276.840000 1419.840000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 267.800000 1419.040000 268.100000 1419.840000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 258.600000 1419.040000 258.900000 1419.840000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 249.860000 1419.040000 250.160000 1419.840000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 241.120000 1419.040000 241.420000 1419.840000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 231.920000 1419.040000 232.220000 1419.840000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 223.180000 1419.040000 223.480000 1419.840000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213.980000 1419.040000 214.280000 1419.840000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.240000 1419.040000 205.540000 1419.840000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.040000 1419.040000 196.340000 1419.840000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 187.300000 1419.040000 187.600000 1419.840000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.560000 1419.040000 178.860000 1419.840000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 169.360000 1419.040000 169.660000 1419.840000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 160.620000 1419.040000 160.920000 1419.840000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 151.420000 1419.040000 151.720000 1419.840000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 142.680000 1419.040000 142.980000 1419.840000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.940000 1419.040000 134.240000 1419.840000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 124.740000 1419.040000 125.040000 1419.840000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.000000 1419.040000 116.300000 1419.840000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 106.800000 1419.040000 107.100000 1419.840000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 98.060000 1419.040000 98.360000 1419.840000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.320000 1419.040000 89.620000 1419.840000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.120000 1419.040000 80.420000 1419.840000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.380000 1419.040000 71.680000 1419.840000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.180000 1419.040000 62.480000 1419.840000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 53.440000 1419.040000 53.740000 1419.840000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.700000 1419.040000 45.000000 1419.840000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 35.500000 1419.040000 35.800000 1419.840000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.760000 1419.040000 27.060000 1419.840000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.560000 1419.040000 17.860000 1419.840000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.820000 1419.040000 9.120000 1419.840000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.080000 1419.040000 0.380000 1419.840000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 651.600000 0.800000 651.900000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 643.060000 0.800000 643.360000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 633.910000 0.800000 634.210000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 625.370000 0.800000 625.670000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 616.220000 0.800000 616.520000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 607.070000 0.800000 607.370000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 598.530000 0.800000 598.830000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 589.380000 0.800000 589.680000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 580.230000 0.800000 580.530000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 571.690000 0.800000 571.990000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 562.540000 0.800000 562.840000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 553.390000 0.800000 553.690000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 544.850000 0.800000 545.150000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 535.700000 0.800000 536.000000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 527.160000 0.800000 527.460000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 518.010000 0.800000 518.310000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 508.860000 0.800000 509.160000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 500.320000 0.800000 500.620000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 491.170000 0.800000 491.470000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 482.020000 0.800000 482.320000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 473.480000 0.800000 473.780000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 464.330000 0.800000 464.630000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 455.790000 0.800000 456.090000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 446.640000 0.800000 446.940000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 437.490000 0.800000 437.790000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 428.950000 0.800000 429.250000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 419.800000 0.800000 420.100000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 410.650000 0.800000 410.950000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 402.110000 0.800000 402.410000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 392.960000 0.800000 393.260000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 384.420000 0.800000 384.720000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 375.270000 0.800000 375.570000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 366.120000 0.800000 366.420000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 357.580000 0.800000 357.880000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 348.430000 0.800000 348.730000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 339.280000 0.800000 339.580000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 330.740000 0.800000 331.040000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 321.590000 0.800000 321.890000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 313.050000 0.800000 313.350000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 303.900000 0.800000 304.200000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 294.750000 0.800000 295.050000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 286.210000 0.800000 286.510000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 277.060000 0.800000 277.360000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 267.910000 0.800000 268.210000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 259.370000 0.800000 259.670000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 250.220000 0.800000 250.520000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 241.070000 0.800000 241.370000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 232.530000 0.800000 232.830000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 223.380000 0.800000 223.680000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 214.840000 0.800000 215.140000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 205.690000 0.800000 205.990000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 196.540000 0.800000 196.840000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 188.000000 0.800000 188.300000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 178.850000 0.800000 179.150000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 169.700000 0.800000 170.000000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 161.160000 0.800000 161.460000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 152.010000 0.800000 152.310000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 143.470000 0.800000 143.770000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 134.320000 0.800000 134.620000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 125.170000 0.800000 125.470000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 116.630000 0.800000 116.930000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 107.480000 0.800000 107.780000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 98.330000 0.800000 98.630000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 89.790000 0.800000 90.090000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 80.640000 0.800000 80.940000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 72.100000 0.800000 72.400000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 62.950000 0.800000 63.250000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 53.800000 0.800000 54.100000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 45.260000 0.800000 45.560000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 36.110000 0.800000 36.410000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 26.960000 0.800000 27.260000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 18.420000 0.800000 18.720000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 9.270000 0.800000 9.570000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1.340000 0.800000 1.640000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1418.370000 0.800000 1418.670000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1410.440000 0.800000 1410.740000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1401.290000 0.800000 1401.590000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1392.750000 0.800000 1393.050000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1383.600000 0.800000 1383.900000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1374.450000 0.800000 1374.750000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1365.910000 0.800000 1366.210000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1356.760000 0.800000 1357.060000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1347.610000 0.800000 1347.910000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1339.070000 0.800000 1339.370000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1329.920000 0.800000 1330.220000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1321.380000 0.800000 1321.680000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1312.230000 0.800000 1312.530000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1303.080000 0.800000 1303.380000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1294.540000 0.800000 1294.840000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1285.390000 0.800000 1285.690000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1276.240000 0.800000 1276.540000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1267.700000 0.800000 1268.000000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1258.550000 0.800000 1258.850000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1250.010000 0.800000 1250.310000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1240.860000 0.800000 1241.160000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1231.710000 0.800000 1232.010000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1223.170000 0.800000 1223.470000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1214.020000 0.800000 1214.320000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1204.870000 0.800000 1205.170000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1196.330000 0.800000 1196.630000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1187.180000 0.800000 1187.480000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1178.640000 0.800000 1178.940000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1169.490000 0.800000 1169.790000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1160.340000 0.800000 1160.640000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1151.800000 0.800000 1152.100000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1142.650000 0.800000 1142.950000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1133.500000 0.800000 1133.800000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1124.960000 0.800000 1125.260000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1115.810000 0.800000 1116.110000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1106.660000 0.800000 1106.960000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1098.120000 0.800000 1098.420000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1088.970000 0.800000 1089.270000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1080.430000 0.800000 1080.730000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1071.280000 0.800000 1071.580000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1062.130000 0.800000 1062.430000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1053.590000 0.800000 1053.890000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1044.440000 0.800000 1044.740000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1035.290000 0.800000 1035.590000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1026.750000 0.800000 1027.050000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1017.600000 0.800000 1017.900000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1009.060000 0.800000 1009.360000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 999.910000 0.800000 1000.210000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 990.760000 0.800000 991.060000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 982.220000 0.800000 982.520000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 973.070000 0.800000 973.370000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 963.920000 0.800000 964.220000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 955.380000 0.800000 955.680000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 946.230000 0.800000 946.530000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 937.690000 0.800000 937.990000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 928.540000 0.800000 928.840000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 919.390000 0.800000 919.690000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 910.850000 0.800000 911.150000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 901.700000 0.800000 902.000000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 892.550000 0.800000 892.850000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 884.010000 0.800000 884.310000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 874.860000 0.800000 875.160000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 866.320000 0.800000 866.620000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 857.170000 0.800000 857.470000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 848.020000 0.800000 848.320000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 839.480000 0.800000 839.780000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 830.330000 0.800000 830.630000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 821.180000 0.800000 821.480000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 812.640000 0.800000 812.940000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 803.490000 0.800000 803.790000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 794.340000 0.800000 794.640000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 785.800000 0.800000 786.100000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 776.650000 0.800000 776.950000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 768.110000 0.800000 768.410000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 758.960000 0.800000 759.260000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 749.810000 0.800000 750.110000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 741.270000 0.800000 741.570000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 732.120000 0.800000 732.420000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 722.970000 0.800000 723.270000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 714.430000 0.800000 714.730000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 705.280000 0.800000 705.580000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 696.740000 0.800000 697.040000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 687.590000 0.800000 687.890000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 678.440000 0.800000 678.740000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 669.900000 0.800000 670.200000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 660.750000 0.800000 661.050000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1053.940000 0.000000 1054.240000 0.800000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1062.680000 0.000000 1062.980000 0.800000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1071.880000 0.000000 1072.180000 0.800000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1080.620000 0.000000 1080.920000 0.800000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1089.360000 0.000000 1089.660000 0.800000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1098.560000 0.000000 1098.860000 0.800000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1107.300000 0.000000 1107.600000 0.800000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1116.500000 0.000000 1116.800000 0.800000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1125.240000 0.000000 1125.540000 0.800000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1133.980000 0.000000 1134.280000 0.800000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1143.180000 0.000000 1143.480000 0.800000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1151.920000 0.000000 1152.220000 0.800000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1161.120000 0.000000 1161.420000 0.800000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1169.860000 0.000000 1170.160000 0.800000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1178.600000 0.000000 1178.900000 0.800000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1187.800000 0.000000 1188.100000 0.800000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.540000 0.000000 1196.840000 0.800000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1205.740000 0.000000 1206.040000 0.800000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1214.480000 0.000000 1214.780000 0.800000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1223.680000 0.000000 1223.980000 0.800000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1232.420000 0.000000 1232.720000 0.800000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1241.160000 0.000000 1241.460000 0.800000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1250.360000 0.000000 1250.660000 0.800000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1259.100000 0.000000 1259.400000 0.800000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1268.300000 0.000000 1268.600000 0.800000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1277.040000 0.000000 1277.340000 0.800000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1285.780000 0.000000 1286.080000 0.800000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1294.980000 0.000000 1295.280000 0.800000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1303.720000 0.000000 1304.020000 0.800000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1312.920000 0.000000 1313.220000 0.800000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1321.660000 0.000000 1321.960000 0.800000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1330.400000 0.000000 1330.700000 0.800000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1339.600000 0.000000 1339.900000 0.800000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1348.340000 0.000000 1348.640000 0.800000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.540000 0.000000 1357.840000 0.800000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1366.280000 0.000000 1366.580000 0.800000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1375.020000 0.000000 1375.320000 0.800000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1384.220000 0.000000 1384.520000 0.800000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1392.960000 0.000000 1393.260000 0.800000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1402.160000 0.000000 1402.460000 0.800000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1410.900000 0.000000 1411.200000 0.800000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.640000 0.000000 1419.940000 0.800000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.080000 0.000000 0.380000 0.800000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 9.280000 0.000000 9.580000 0.800000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.020000 0.000000 18.320000 0.800000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 27.220000 0.000000 27.520000 0.800000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 35.960000 0.000000 36.260000 0.800000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.160000 0.000000 45.460000 0.800000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 53.900000 0.000000 54.200000 0.800000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.640000 0.000000 62.940000 0.800000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.840000 0.000000 72.140000 0.800000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.580000 0.000000 80.880000 0.800000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.780000 0.000000 90.080000 0.800000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 98.520000 0.000000 98.820000 0.800000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.260000 0.000000 107.560000 0.800000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.460000 0.000000 116.760000 0.800000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 125.200000 0.000000 125.500000 0.800000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 134.400000 0.000000 134.700000 0.800000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 143.140000 0.000000 143.440000 0.800000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 151.880000 0.000000 152.180000 0.800000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.080000 0.000000 161.380000 0.800000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 169.820000 0.000000 170.120000 0.800000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 179.020000 0.000000 179.320000 0.800000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 187.760000 0.000000 188.060000 0.800000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.500000 0.000000 196.800000 0.800000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.700000 0.000000 206.000000 0.800000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 214.440000 0.000000 214.740000 0.800000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 223.640000 0.000000 223.940000 0.800000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.380000 0.000000 232.680000 0.800000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 241.580000 0.000000 241.880000 0.800000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.320000 0.000000 250.620000 0.800000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 259.060000 0.000000 259.360000 0.800000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.260000 0.000000 268.560000 0.800000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 277.000000 0.000000 277.300000 0.800000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 286.200000 0.000000 286.500000 0.800000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 294.940000 0.000000 295.240000 0.800000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 303.680000 0.000000 303.980000 0.800000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 312.880000 0.000000 313.180000 0.800000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 321.620000 0.000000 321.920000 0.800000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 330.820000 0.000000 331.120000 0.800000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 339.560000 0.000000 339.860000 0.800000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 348.300000 0.000000 348.600000 0.800000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 357.500000 0.000000 357.800000 0.800000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 366.240000 0.000000 366.540000 0.800000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 375.440000 0.000000 375.740000 0.800000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 384.180000 0.000000 384.480000 0.800000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 392.920000 0.000000 393.220000 0.800000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 402.120000 0.000000 402.420000 0.800000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 410.860000 0.000000 411.160000 0.800000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 420.060000 0.000000 420.360000 0.800000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 428.800000 0.000000 429.100000 0.800000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 438.000000 0.000000 438.300000 0.800000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.740000 0.000000 447.040000 0.800000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 455.480000 0.000000 455.780000 0.800000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 464.680000 0.000000 464.980000 0.800000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.420000 0.000000 473.720000 0.800000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 482.620000 0.000000 482.920000 0.800000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 491.360000 0.000000 491.660000 0.800000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.100000 0.000000 500.400000 0.800000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 509.300000 0.000000 509.600000 0.800000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 518.040000 0.000000 518.340000 0.800000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 527.240000 0.000000 527.540000 0.800000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 535.980000 0.000000 536.280000 0.800000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 544.720000 0.000000 545.020000 0.800000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 553.920000 0.000000 554.220000 0.800000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 562.660000 0.000000 562.960000 0.800000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 571.860000 0.000000 572.160000 0.800000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 580.600000 0.000000 580.900000 0.800000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 589.340000 0.000000 589.640000 0.800000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 598.540000 0.000000 598.840000 0.800000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 607.280000 0.000000 607.580000 0.800000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 616.480000 0.000000 616.780000 0.800000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 625.220000 0.000000 625.520000 0.800000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 634.420000 0.000000 634.720000 0.800000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 643.160000 0.000000 643.460000 0.800000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 651.900000 0.000000 652.200000 0.800000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 661.100000 0.000000 661.400000 0.800000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 669.840000 0.000000 670.140000 0.800000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 679.040000 0.000000 679.340000 0.800000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 687.780000 0.000000 688.080000 0.800000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.520000 0.000000 696.820000 0.800000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 705.720000 0.000000 706.020000 0.800000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 714.460000 0.000000 714.760000 0.800000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 723.660000 0.000000 723.960000 0.800000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 732.400000 0.000000 732.700000 0.800000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 741.140000 0.000000 741.440000 0.800000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 750.340000 0.000000 750.640000 0.800000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 759.080000 0.000000 759.380000 0.800000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 768.280000 0.000000 768.580000 0.800000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 777.020000 0.000000 777.320000 0.800000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 785.760000 0.000000 786.060000 0.800000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 794.960000 0.000000 795.260000 0.800000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 803.700000 0.000000 804.000000 0.800000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 812.900000 0.000000 813.200000 0.800000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 821.640000 0.000000 821.940000 0.800000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 830.840000 0.000000 831.140000 0.800000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 839.580000 0.000000 839.880000 0.800000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 848.320000 0.000000 848.620000 0.800000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 857.520000 0.000000 857.820000 0.800000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 866.260000 0.000000 866.560000 0.800000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 875.460000 0.000000 875.760000 0.800000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 884.200000 0.000000 884.500000 0.800000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 892.940000 0.000000 893.240000 0.800000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 902.140000 0.000000 902.440000 0.800000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 910.880000 0.000000 911.180000 0.800000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 920.080000 0.000000 920.380000 0.800000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.820000 0.000000 929.120000 0.800000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 937.560000 0.000000 937.860000 0.800000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 946.760000 0.000000 947.060000 0.800000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 955.500000 0.000000 955.800000 0.800000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 964.700000 0.000000 965.000000 0.800000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 973.440000 0.000000 973.740000 0.800000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 982.180000 0.000000 982.480000 0.800000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 991.380000 0.000000 991.680000 0.800000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1000.120000 0.000000 1000.420000 0.800000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1009.320000 0.000000 1009.620000 0.800000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1018.060000 0.000000 1018.360000 0.800000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1027.260000 0.000000 1027.560000 0.800000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1036.000000 0.000000 1036.300000 0.800000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1044.740000 0.000000 1045.040000 0.800000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 37.330000 1420.020000 37.630000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 46.480000 1420.020000 46.780000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 55.630000 1420.020000 55.930000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 64.780000 1420.020000 65.080000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 73.930000 1420.020000 74.230000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 83.080000 1420.020000 83.380000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 92.230000 1420.020000 92.530000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 101.380000 1420.020000 101.680000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 109.920000 1420.020000 110.220000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 119.070000 1420.020000 119.370000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 819.350000 1420.020000 819.650000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 828.500000 1420.020000 828.800000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 837.650000 1420.020000 837.950000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 846.800000 1420.020000 847.100000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 855.950000 1420.020000 856.250000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 865.100000 1420.020000 865.400000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 874.250000 1420.020000 874.550000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 883.400000 1420.020000 883.700000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 892.550000 1420.020000 892.850000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 901.700000 1420.020000 902.000000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 910.850000 1420.020000 911.150000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 919.390000 1420.020000 919.690000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 928.540000 1420.020000 928.840000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 937.690000 1420.020000 937.990000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 946.840000 1420.020000 947.140000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 955.990000 1420.020000 956.290000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 965.140000 1420.020000 965.440000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 974.290000 1420.020000 974.590000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 983.440000 1420.020000 983.740000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 992.590000 1420.020000 992.890000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1001.740000 1420.020000 1002.040000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1010.890000 1420.020000 1011.190000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1019.430000 1420.020000 1019.730000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1028.580000 1420.020000 1028.880000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1037.730000 1420.020000 1038.030000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1046.880000 1420.020000 1047.180000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1056.030000 1420.020000 1056.330000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1065.180000 1420.020000 1065.480000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1074.330000 1420.020000 1074.630000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1083.480000 1420.020000 1083.780000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1092.630000 1420.020000 1092.930000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1101.780000 1420.020000 1102.080000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1110.930000 1420.020000 1111.230000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1119.470000 1420.020000 1119.770000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1128.620000 1420.020000 1128.920000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1137.770000 1420.020000 1138.070000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1146.920000 1420.020000 1147.220000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1156.070000 1420.020000 1156.370000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 128.220000 1420.020000 128.520000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 137.370000 1420.020000 137.670000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 146.520000 1420.020000 146.820000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 155.670000 1420.020000 155.970000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 164.820000 1420.020000 165.120000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 173.970000 1420.020000 174.270000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 183.120000 1420.020000 183.420000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 192.270000 1420.020000 192.570000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 201.420000 1420.020000 201.720000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 209.960000 1420.020000 210.260000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 219.110000 1420.020000 219.410000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 228.260000 1420.020000 228.560000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 237.410000 1420.020000 237.710000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 246.560000 1420.020000 246.860000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 255.710000 1420.020000 256.010000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 264.860000 1420.020000 265.160000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 274.010000 1420.020000 274.310000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 283.160000 1420.020000 283.460000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 292.310000 1420.020000 292.610000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 301.460000 1420.020000 301.760000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 310.000000 1420.020000 310.300000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 319.150000 1420.020000 319.450000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 328.300000 1420.020000 328.600000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 337.450000 1420.020000 337.750000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 346.600000 1420.020000 346.900000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 355.750000 1420.020000 356.050000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 364.900000 1420.020000 365.200000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 374.050000 1420.020000 374.350000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 383.200000 1420.020000 383.500000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 392.350000 1420.020000 392.650000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 401.500000 1420.020000 401.800000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 410.040000 1420.020000 410.340000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 419.190000 1420.020000 419.490000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 428.340000 1420.020000 428.640000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 437.490000 1420.020000 437.790000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 446.640000 1420.020000 446.940000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 455.790000 1420.020000 456.090000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 464.940000 1420.020000 465.240000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 474.090000 1420.020000 474.390000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 483.240000 1420.020000 483.540000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 492.390000 1420.020000 492.690000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 501.540000 1420.020000 501.840000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 510.080000 1420.020000 510.380000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 519.230000 1420.020000 519.530000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 528.380000 1420.020000 528.680000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 537.530000 1420.020000 537.830000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 546.680000 1420.020000 546.980000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 555.830000 1420.020000 556.130000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 564.980000 1420.020000 565.280000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 574.130000 1420.020000 574.430000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 583.280000 1420.020000 583.580000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 592.430000 1420.020000 592.730000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 601.580000 1420.020000 601.880000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 610.120000 1420.020000 610.420000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 619.270000 1420.020000 619.570000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 628.420000 1420.020000 628.720000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 637.570000 1420.020000 637.870000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 646.720000 1420.020000 647.020000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 655.870000 1420.020000 656.170000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 665.020000 1420.020000 665.320000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 674.170000 1420.020000 674.470000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 683.320000 1420.020000 683.620000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 692.470000 1420.020000 692.770000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 701.620000 1420.020000 701.920000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 710.160000 1420.020000 710.460000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 719.310000 1420.020000 719.610000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 728.460000 1420.020000 728.760000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 737.610000 1420.020000 737.910000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 746.760000 1420.020000 747.060000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 755.910000 1420.020000 756.210000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 765.060000 1420.020000 765.360000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 774.210000 1420.020000 774.510000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 783.360000 1420.020000 783.660000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 792.510000 1420.020000 792.810000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 801.660000 1420.020000 801.960000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 810.810000 1420.020000 811.110000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1165.220000 1420.020000 1165.520000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1174.370000 1420.020000 1174.670000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1183.520000 1420.020000 1183.820000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1192.670000 1420.020000 1192.970000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1201.820000 1420.020000 1202.120000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1210.970000 1420.020000 1211.270000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1219.510000 1420.020000 1219.810000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1228.660000 1420.020000 1228.960000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1237.810000 1420.020000 1238.110000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1246.960000 1420.020000 1247.260000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1256.110000 1420.020000 1256.410000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1265.260000 1420.020000 1265.560000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1274.410000 1420.020000 1274.710000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1283.560000 1420.020000 1283.860000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1292.710000 1420.020000 1293.010000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1301.860000 1420.020000 1302.160000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1311.010000 1420.020000 1311.310000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1319.550000 1420.020000 1319.850000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1328.700000 1420.020000 1329.000000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1337.850000 1420.020000 1338.150000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1347.000000 1420.020000 1347.300000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1356.150000 1420.020000 1356.450000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1365.300000 1420.020000 1365.600000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1374.450000 1420.020000 1374.750000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1383.600000 1420.020000 1383.900000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1392.750000 1420.020000 1393.050000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1401.900000 1420.020000 1402.200000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1411.050000 1420.020000 1411.350000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1418.370000 1420.020000 1418.670000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 28.180000 1420.020000 28.480000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 1.340000 1420.020000 1.640000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 9.880000 1420.020000 10.180000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1419.220000 19.030000 1420.020000 19.330000 ;
    END
  END user_irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 2.520000 2.260000 1417.500000 4.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.520000 1413.540000 1417.500000 1415.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1415.500000 2.260000 1417.500000 1415.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.520000 2.260000 4.520000 1415.540000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.520000 2.260000 4.520000 1415.540000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1195.325000 811.465000 1197.065000 1206.245000 ;
      LAYER met4 ;
        RECT 720.005000 811.465000 721.745000 1206.245000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 681.545000 811.465000 683.285000 1206.245000 ;
      LAYER met4 ;
        RECT 206.225000 811.465000 207.965000 1206.245000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 6.320000 6.060000 1413.700000 8.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.320000 1409.740000 1413.700000 1411.740000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1411.700000 6.060000 1413.700000 1411.740000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.320000 6.060000 8.320000 1411.740000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 723.405000 814.865000 725.145000 1202.845000 ;
      LAYER met4 ;
        RECT 1191.925000 814.865000 1193.665000 1202.845000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 209.625000 814.865000 211.365000 1202.845000 ;
      LAYER met4 ;
        RECT 678.145000 814.865000 679.885000 1202.845000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 1415.710000 1420.020000 1419.840000 ;
      RECT 4.690000 2.090000 1420.020000 1415.710000 ;
      RECT 0.000000 2.090000 2.350000 1415.710000 ;
      RECT 0.000000 0.000000 1420.020000 2.090000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1420.020000 1419.840000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 1420.020000 1419.840000 ;
    LAYER met3 ;
      RECT 1411.040000 1418.970000 1419.340000 1419.840000 ;
      RECT 0.680000 1418.970000 8.520000 1419.840000 ;
      RECT 1411.040000 1418.740000 1418.920000 1418.970000 ;
      RECT 1402.300000 1418.740000 1410.140000 1419.840000 ;
      RECT 1393.100000 1418.740000 1401.400000 1419.840000 ;
      RECT 1384.360000 1418.740000 1392.200000 1419.840000 ;
      RECT 1375.160000 1418.740000 1383.460000 1419.840000 ;
      RECT 1366.420000 1418.740000 1374.260000 1419.840000 ;
      RECT 1357.680000 1418.740000 1365.520000 1419.840000 ;
      RECT 1348.480000 1418.740000 1356.780000 1419.840000 ;
      RECT 1339.740000 1418.740000 1347.580000 1419.840000 ;
      RECT 1330.540000 1418.740000 1338.840000 1419.840000 ;
      RECT 1321.800000 1418.740000 1329.640000 1419.840000 ;
      RECT 1313.060000 1418.740000 1320.900000 1419.840000 ;
      RECT 1303.860000 1418.740000 1312.160000 1419.840000 ;
      RECT 1295.120000 1418.740000 1302.960000 1419.840000 ;
      RECT 1285.920000 1418.740000 1294.220000 1419.840000 ;
      RECT 1277.180000 1418.740000 1285.020000 1419.840000 ;
      RECT 1268.440000 1418.740000 1276.280000 1419.840000 ;
      RECT 1259.240000 1418.740000 1267.540000 1419.840000 ;
      RECT 1250.500000 1418.740000 1258.340000 1419.840000 ;
      RECT 1241.300000 1418.740000 1249.600000 1419.840000 ;
      RECT 1232.560000 1418.740000 1240.400000 1419.840000 ;
      RECT 1223.820000 1418.740000 1231.660000 1419.840000 ;
      RECT 1214.620000 1418.740000 1222.920000 1419.840000 ;
      RECT 1205.880000 1418.740000 1213.720000 1419.840000 ;
      RECT 1196.680000 1418.740000 1204.980000 1419.840000 ;
      RECT 1187.940000 1418.740000 1195.780000 1419.840000 ;
      RECT 1178.740000 1418.740000 1187.040000 1419.840000 ;
      RECT 1170.000000 1418.740000 1177.840000 1419.840000 ;
      RECT 1161.260000 1418.740000 1169.100000 1419.840000 ;
      RECT 1152.060000 1418.740000 1160.360000 1419.840000 ;
      RECT 1143.320000 1418.740000 1151.160000 1419.840000 ;
      RECT 1134.120000 1418.740000 1142.420000 1419.840000 ;
      RECT 1125.380000 1418.740000 1133.220000 1419.840000 ;
      RECT 1116.640000 1418.740000 1124.480000 1419.840000 ;
      RECT 1107.440000 1418.740000 1115.740000 1419.840000 ;
      RECT 1098.700000 1418.740000 1106.540000 1419.840000 ;
      RECT 1089.500000 1418.740000 1097.800000 1419.840000 ;
      RECT 1080.760000 1418.740000 1088.600000 1419.840000 ;
      RECT 1072.020000 1418.740000 1079.860000 1419.840000 ;
      RECT 1062.820000 1418.740000 1071.120000 1419.840000 ;
      RECT 1054.080000 1418.740000 1061.920000 1419.840000 ;
      RECT 1044.880000 1418.740000 1053.180000 1419.840000 ;
      RECT 1036.140000 1418.740000 1043.980000 1419.840000 ;
      RECT 1027.400000 1418.740000 1035.240000 1419.840000 ;
      RECT 1018.200000 1418.740000 1026.500000 1419.840000 ;
      RECT 1009.460000 1418.740000 1017.300000 1419.840000 ;
      RECT 1000.260000 1418.740000 1008.560000 1419.840000 ;
      RECT 991.520000 1418.740000 999.360000 1419.840000 ;
      RECT 982.320000 1418.740000 990.620000 1419.840000 ;
      RECT 973.580000 1418.740000 981.420000 1419.840000 ;
      RECT 964.840000 1418.740000 972.680000 1419.840000 ;
      RECT 955.640000 1418.740000 963.940000 1419.840000 ;
      RECT 946.900000 1418.740000 954.740000 1419.840000 ;
      RECT 937.700000 1418.740000 946.000000 1419.840000 ;
      RECT 928.960000 1418.740000 936.800000 1419.840000 ;
      RECT 920.220000 1418.740000 928.060000 1419.840000 ;
      RECT 911.020000 1418.740000 919.320000 1419.840000 ;
      RECT 902.280000 1418.740000 910.120000 1419.840000 ;
      RECT 893.080000 1418.740000 901.380000 1419.840000 ;
      RECT 884.340000 1418.740000 892.180000 1419.840000 ;
      RECT 875.600000 1418.740000 883.440000 1419.840000 ;
      RECT 866.400000 1418.740000 874.700000 1419.840000 ;
      RECT 857.660000 1418.740000 865.500000 1419.840000 ;
      RECT 848.460000 1418.740000 856.760000 1419.840000 ;
      RECT 839.720000 1418.740000 847.560000 1419.840000 ;
      RECT 830.980000 1418.740000 838.820000 1419.840000 ;
      RECT 821.780000 1418.740000 830.080000 1419.840000 ;
      RECT 813.040000 1418.740000 820.880000 1419.840000 ;
      RECT 803.840000 1418.740000 812.140000 1419.840000 ;
      RECT 795.100000 1418.740000 802.940000 1419.840000 ;
      RECT 785.900000 1418.740000 794.200000 1419.840000 ;
      RECT 777.160000 1418.740000 785.000000 1419.840000 ;
      RECT 768.420000 1418.740000 776.260000 1419.840000 ;
      RECT 759.220000 1418.740000 767.520000 1419.840000 ;
      RECT 750.480000 1418.740000 758.320000 1419.840000 ;
      RECT 741.280000 1418.740000 749.580000 1419.840000 ;
      RECT 732.540000 1418.740000 740.380000 1419.840000 ;
      RECT 723.800000 1418.740000 731.640000 1419.840000 ;
      RECT 714.600000 1418.740000 722.900000 1419.840000 ;
      RECT 705.860000 1418.740000 713.700000 1419.840000 ;
      RECT 696.660000 1418.740000 704.960000 1419.840000 ;
      RECT 687.920000 1418.740000 695.760000 1419.840000 ;
      RECT 679.180000 1418.740000 687.020000 1419.840000 ;
      RECT 669.980000 1418.740000 678.280000 1419.840000 ;
      RECT 661.240000 1418.740000 669.080000 1419.840000 ;
      RECT 652.040000 1418.740000 660.340000 1419.840000 ;
      RECT 643.300000 1418.740000 651.140000 1419.840000 ;
      RECT 634.560000 1418.740000 642.400000 1419.840000 ;
      RECT 625.360000 1418.740000 633.660000 1419.840000 ;
      RECT 616.620000 1418.740000 624.460000 1419.840000 ;
      RECT 607.420000 1418.740000 615.720000 1419.840000 ;
      RECT 598.680000 1418.740000 606.520000 1419.840000 ;
      RECT 589.480000 1418.740000 597.780000 1419.840000 ;
      RECT 580.740000 1418.740000 588.580000 1419.840000 ;
      RECT 572.000000 1418.740000 579.840000 1419.840000 ;
      RECT 562.800000 1418.740000 571.100000 1419.840000 ;
      RECT 554.060000 1418.740000 561.900000 1419.840000 ;
      RECT 544.860000 1418.740000 553.160000 1419.840000 ;
      RECT 536.120000 1418.740000 543.960000 1419.840000 ;
      RECT 527.380000 1418.740000 535.220000 1419.840000 ;
      RECT 518.180000 1418.740000 526.480000 1419.840000 ;
      RECT 509.440000 1418.740000 517.280000 1419.840000 ;
      RECT 500.240000 1418.740000 508.540000 1419.840000 ;
      RECT 491.500000 1418.740000 499.340000 1419.840000 ;
      RECT 482.760000 1418.740000 490.600000 1419.840000 ;
      RECT 473.560000 1418.740000 481.860000 1419.840000 ;
      RECT 464.820000 1418.740000 472.660000 1419.840000 ;
      RECT 455.620000 1418.740000 463.920000 1419.840000 ;
      RECT 446.880000 1418.740000 454.720000 1419.840000 ;
      RECT 438.140000 1418.740000 445.980000 1419.840000 ;
      RECT 428.940000 1418.740000 437.240000 1419.840000 ;
      RECT 420.200000 1418.740000 428.040000 1419.840000 ;
      RECT 411.000000 1418.740000 419.300000 1419.840000 ;
      RECT 402.260000 1418.740000 410.100000 1419.840000 ;
      RECT 393.060000 1418.740000 401.360000 1419.840000 ;
      RECT 384.320000 1418.740000 392.160000 1419.840000 ;
      RECT 375.580000 1418.740000 383.420000 1419.840000 ;
      RECT 366.380000 1418.740000 374.680000 1419.840000 ;
      RECT 357.640000 1418.740000 365.480000 1419.840000 ;
      RECT 348.440000 1418.740000 356.740000 1419.840000 ;
      RECT 339.700000 1418.740000 347.540000 1419.840000 ;
      RECT 330.960000 1418.740000 338.800000 1419.840000 ;
      RECT 321.760000 1418.740000 330.060000 1419.840000 ;
      RECT 313.020000 1418.740000 320.860000 1419.840000 ;
      RECT 303.820000 1418.740000 312.120000 1419.840000 ;
      RECT 295.080000 1418.740000 302.920000 1419.840000 ;
      RECT 286.340000 1418.740000 294.180000 1419.840000 ;
      RECT 277.140000 1418.740000 285.440000 1419.840000 ;
      RECT 268.400000 1418.740000 276.240000 1419.840000 ;
      RECT 259.200000 1418.740000 267.500000 1419.840000 ;
      RECT 250.460000 1418.740000 258.300000 1419.840000 ;
      RECT 241.720000 1418.740000 249.560000 1419.840000 ;
      RECT 232.520000 1418.740000 240.820000 1419.840000 ;
      RECT 223.780000 1418.740000 231.620000 1419.840000 ;
      RECT 214.580000 1418.740000 222.880000 1419.840000 ;
      RECT 205.840000 1418.740000 213.680000 1419.840000 ;
      RECT 196.640000 1418.740000 204.940000 1419.840000 ;
      RECT 187.900000 1418.740000 195.740000 1419.840000 ;
      RECT 179.160000 1418.740000 187.000000 1419.840000 ;
      RECT 169.960000 1418.740000 178.260000 1419.840000 ;
      RECT 161.220000 1418.740000 169.060000 1419.840000 ;
      RECT 152.020000 1418.740000 160.320000 1419.840000 ;
      RECT 143.280000 1418.740000 151.120000 1419.840000 ;
      RECT 134.540000 1418.740000 142.380000 1419.840000 ;
      RECT 125.340000 1418.740000 133.640000 1419.840000 ;
      RECT 116.600000 1418.740000 124.440000 1419.840000 ;
      RECT 107.400000 1418.740000 115.700000 1419.840000 ;
      RECT 98.660000 1418.740000 106.500000 1419.840000 ;
      RECT 89.920000 1418.740000 97.760000 1419.840000 ;
      RECT 80.720000 1418.740000 89.020000 1419.840000 ;
      RECT 71.980000 1418.740000 79.820000 1419.840000 ;
      RECT 62.780000 1418.740000 71.080000 1419.840000 ;
      RECT 54.040000 1418.740000 61.880000 1419.840000 ;
      RECT 45.300000 1418.740000 53.140000 1419.840000 ;
      RECT 36.100000 1418.740000 44.400000 1419.840000 ;
      RECT 27.360000 1418.740000 35.200000 1419.840000 ;
      RECT 18.160000 1418.740000 26.460000 1419.840000 ;
      RECT 9.420000 1418.740000 17.260000 1419.840000 ;
      RECT 1.100000 1418.740000 8.520000 1418.970000 ;
      RECT 1.100000 1418.070000 1418.920000 1418.740000 ;
      RECT 0.000000 1415.840000 1420.020000 1418.070000 ;
      RECT 1417.800000 1413.240000 1420.020000 1415.840000 ;
      RECT 0.000000 1413.240000 2.220000 1415.840000 ;
      RECT 0.000000 1412.040000 1420.020000 1413.240000 ;
      RECT 1414.000000 1411.650000 1420.020000 1412.040000 ;
      RECT 0.000000 1411.040000 6.020000 1412.040000 ;
      RECT 1414.000000 1410.750000 1418.920000 1411.650000 ;
      RECT 1.100000 1410.140000 6.020000 1411.040000 ;
      RECT 1414.000000 1409.440000 1420.020000 1410.750000 ;
      RECT 0.000000 1409.440000 6.020000 1410.140000 ;
      RECT 0.000000 1402.500000 1420.020000 1409.440000 ;
      RECT 0.000000 1401.890000 1418.920000 1402.500000 ;
      RECT 1.100000 1401.600000 1418.920000 1401.890000 ;
      RECT 1.100000 1400.990000 1420.020000 1401.600000 ;
      RECT 0.000000 1393.350000 1420.020000 1400.990000 ;
      RECT 1.100000 1392.450000 1418.920000 1393.350000 ;
      RECT 0.000000 1384.200000 1420.020000 1392.450000 ;
      RECT 1.100000 1383.300000 1418.920000 1384.200000 ;
      RECT 0.000000 1375.050000 1420.020000 1383.300000 ;
      RECT 1.100000 1374.150000 1418.920000 1375.050000 ;
      RECT 0.000000 1366.510000 1420.020000 1374.150000 ;
      RECT 1.100000 1365.900000 1420.020000 1366.510000 ;
      RECT 1.100000 1365.610000 1418.920000 1365.900000 ;
      RECT 0.000000 1365.000000 1418.920000 1365.610000 ;
      RECT 0.000000 1357.360000 1420.020000 1365.000000 ;
      RECT 1.100000 1356.750000 1420.020000 1357.360000 ;
      RECT 1.100000 1356.460000 1418.920000 1356.750000 ;
      RECT 0.000000 1355.850000 1418.920000 1356.460000 ;
      RECT 0.000000 1348.210000 1420.020000 1355.850000 ;
      RECT 1.100000 1347.600000 1420.020000 1348.210000 ;
      RECT 1.100000 1347.310000 1418.920000 1347.600000 ;
      RECT 0.000000 1346.700000 1418.920000 1347.310000 ;
      RECT 0.000000 1339.670000 1420.020000 1346.700000 ;
      RECT 1.100000 1338.770000 1420.020000 1339.670000 ;
      RECT 0.000000 1338.450000 1420.020000 1338.770000 ;
      RECT 0.000000 1337.550000 1418.920000 1338.450000 ;
      RECT 0.000000 1330.520000 1420.020000 1337.550000 ;
      RECT 1.100000 1329.620000 1420.020000 1330.520000 ;
      RECT 0.000000 1329.300000 1420.020000 1329.620000 ;
      RECT 0.000000 1328.400000 1418.920000 1329.300000 ;
      RECT 0.000000 1321.980000 1420.020000 1328.400000 ;
      RECT 1.100000 1321.080000 1420.020000 1321.980000 ;
      RECT 0.000000 1320.150000 1420.020000 1321.080000 ;
      RECT 0.000000 1319.250000 1418.920000 1320.150000 ;
      RECT 0.000000 1312.830000 1420.020000 1319.250000 ;
      RECT 1.100000 1311.930000 1420.020000 1312.830000 ;
      RECT 0.000000 1311.610000 1420.020000 1311.930000 ;
      RECT 0.000000 1310.710000 1418.920000 1311.610000 ;
      RECT 0.000000 1303.680000 1420.020000 1310.710000 ;
      RECT 1.100000 1302.780000 1420.020000 1303.680000 ;
      RECT 0.000000 1302.460000 1420.020000 1302.780000 ;
      RECT 0.000000 1301.560000 1418.920000 1302.460000 ;
      RECT 0.000000 1295.140000 1420.020000 1301.560000 ;
      RECT 1.100000 1294.240000 1420.020000 1295.140000 ;
      RECT 0.000000 1293.310000 1420.020000 1294.240000 ;
      RECT 0.000000 1292.410000 1418.920000 1293.310000 ;
      RECT 0.000000 1285.990000 1420.020000 1292.410000 ;
      RECT 1.100000 1285.090000 1420.020000 1285.990000 ;
      RECT 0.000000 1284.160000 1420.020000 1285.090000 ;
      RECT 0.000000 1283.260000 1418.920000 1284.160000 ;
      RECT 0.000000 1276.840000 1420.020000 1283.260000 ;
      RECT 1.100000 1275.940000 1420.020000 1276.840000 ;
      RECT 0.000000 1275.010000 1420.020000 1275.940000 ;
      RECT 0.000000 1274.110000 1418.920000 1275.010000 ;
      RECT 0.000000 1268.300000 1420.020000 1274.110000 ;
      RECT 1.100000 1267.400000 1420.020000 1268.300000 ;
      RECT 0.000000 1265.860000 1420.020000 1267.400000 ;
      RECT 0.000000 1264.960000 1418.920000 1265.860000 ;
      RECT 0.000000 1259.150000 1420.020000 1264.960000 ;
      RECT 1.100000 1258.250000 1420.020000 1259.150000 ;
      RECT 0.000000 1256.710000 1420.020000 1258.250000 ;
      RECT 0.000000 1255.810000 1418.920000 1256.710000 ;
      RECT 0.000000 1250.610000 1420.020000 1255.810000 ;
      RECT 1.100000 1249.710000 1420.020000 1250.610000 ;
      RECT 0.000000 1247.560000 1420.020000 1249.710000 ;
      RECT 0.000000 1246.660000 1418.920000 1247.560000 ;
      RECT 0.000000 1241.460000 1420.020000 1246.660000 ;
      RECT 1.100000 1240.560000 1420.020000 1241.460000 ;
      RECT 0.000000 1238.410000 1420.020000 1240.560000 ;
      RECT 0.000000 1237.510000 1418.920000 1238.410000 ;
      RECT 0.000000 1232.310000 1420.020000 1237.510000 ;
      RECT 1.100000 1231.410000 1420.020000 1232.310000 ;
      RECT 0.000000 1229.260000 1420.020000 1231.410000 ;
      RECT 0.000000 1228.360000 1418.920000 1229.260000 ;
      RECT 0.000000 1223.770000 1420.020000 1228.360000 ;
      RECT 1.100000 1222.870000 1420.020000 1223.770000 ;
      RECT 0.000000 1220.110000 1420.020000 1222.870000 ;
      RECT 0.000000 1219.210000 1418.920000 1220.110000 ;
      RECT 0.000000 1214.620000 1420.020000 1219.210000 ;
      RECT 1.100000 1213.720000 1420.020000 1214.620000 ;
      RECT 0.000000 1211.570000 1420.020000 1213.720000 ;
      RECT 0.000000 1210.670000 1418.920000 1211.570000 ;
      RECT 0.000000 1205.470000 1420.020000 1210.670000 ;
      RECT 1.100000 1204.570000 1420.020000 1205.470000 ;
      RECT 0.000000 1202.420000 1420.020000 1204.570000 ;
      RECT 0.000000 1201.520000 1418.920000 1202.420000 ;
      RECT 0.000000 1196.930000 1420.020000 1201.520000 ;
      RECT 1.100000 1196.030000 1420.020000 1196.930000 ;
      RECT 0.000000 1193.270000 1420.020000 1196.030000 ;
      RECT 0.000000 1192.370000 1418.920000 1193.270000 ;
      RECT 0.000000 1187.780000 1420.020000 1192.370000 ;
      RECT 1.100000 1186.880000 1420.020000 1187.780000 ;
      RECT 0.000000 1184.120000 1420.020000 1186.880000 ;
      RECT 0.000000 1183.220000 1418.920000 1184.120000 ;
      RECT 0.000000 1179.240000 1420.020000 1183.220000 ;
      RECT 1.100000 1178.340000 1420.020000 1179.240000 ;
      RECT 0.000000 1174.970000 1420.020000 1178.340000 ;
      RECT 0.000000 1174.070000 1418.920000 1174.970000 ;
      RECT 0.000000 1170.090000 1420.020000 1174.070000 ;
      RECT 1.100000 1169.190000 1420.020000 1170.090000 ;
      RECT 0.000000 1165.820000 1420.020000 1169.190000 ;
      RECT 0.000000 1164.920000 1418.920000 1165.820000 ;
      RECT 0.000000 1160.940000 1420.020000 1164.920000 ;
      RECT 1.100000 1160.040000 1420.020000 1160.940000 ;
      RECT 0.000000 1156.670000 1420.020000 1160.040000 ;
      RECT 0.000000 1155.770000 1418.920000 1156.670000 ;
      RECT 0.000000 1152.400000 1420.020000 1155.770000 ;
      RECT 1.100000 1151.500000 1420.020000 1152.400000 ;
      RECT 0.000000 1147.520000 1420.020000 1151.500000 ;
      RECT 0.000000 1146.620000 1418.920000 1147.520000 ;
      RECT 0.000000 1143.250000 1420.020000 1146.620000 ;
      RECT 1.100000 1142.350000 1420.020000 1143.250000 ;
      RECT 0.000000 1138.370000 1420.020000 1142.350000 ;
      RECT 0.000000 1137.470000 1418.920000 1138.370000 ;
      RECT 0.000000 1134.100000 1420.020000 1137.470000 ;
      RECT 1.100000 1133.200000 1420.020000 1134.100000 ;
      RECT 0.000000 1129.220000 1420.020000 1133.200000 ;
      RECT 0.000000 1128.320000 1418.920000 1129.220000 ;
      RECT 0.000000 1125.560000 1420.020000 1128.320000 ;
      RECT 1.100000 1124.660000 1420.020000 1125.560000 ;
      RECT 0.000000 1120.070000 1420.020000 1124.660000 ;
      RECT 0.000000 1119.170000 1418.920000 1120.070000 ;
      RECT 0.000000 1116.410000 1420.020000 1119.170000 ;
      RECT 1.100000 1115.510000 1420.020000 1116.410000 ;
      RECT 0.000000 1111.530000 1420.020000 1115.510000 ;
      RECT 0.000000 1110.630000 1418.920000 1111.530000 ;
      RECT 0.000000 1107.260000 1420.020000 1110.630000 ;
      RECT 1.100000 1106.360000 1420.020000 1107.260000 ;
      RECT 0.000000 1102.380000 1420.020000 1106.360000 ;
      RECT 0.000000 1101.480000 1418.920000 1102.380000 ;
      RECT 0.000000 1098.720000 1420.020000 1101.480000 ;
      RECT 1.100000 1097.820000 1420.020000 1098.720000 ;
      RECT 0.000000 1093.230000 1420.020000 1097.820000 ;
      RECT 0.000000 1092.330000 1418.920000 1093.230000 ;
      RECT 0.000000 1089.570000 1420.020000 1092.330000 ;
      RECT 1.100000 1088.670000 1420.020000 1089.570000 ;
      RECT 0.000000 1084.080000 1420.020000 1088.670000 ;
      RECT 0.000000 1083.180000 1418.920000 1084.080000 ;
      RECT 0.000000 1081.030000 1420.020000 1083.180000 ;
      RECT 1.100000 1080.130000 1420.020000 1081.030000 ;
      RECT 0.000000 1074.930000 1420.020000 1080.130000 ;
      RECT 0.000000 1074.030000 1418.920000 1074.930000 ;
      RECT 0.000000 1071.880000 1420.020000 1074.030000 ;
      RECT 1.100000 1070.980000 1420.020000 1071.880000 ;
      RECT 0.000000 1065.780000 1420.020000 1070.980000 ;
      RECT 0.000000 1064.880000 1418.920000 1065.780000 ;
      RECT 0.000000 1062.730000 1420.020000 1064.880000 ;
      RECT 1.100000 1061.830000 1420.020000 1062.730000 ;
      RECT 0.000000 1056.630000 1420.020000 1061.830000 ;
      RECT 0.000000 1055.730000 1418.920000 1056.630000 ;
      RECT 0.000000 1054.190000 1420.020000 1055.730000 ;
      RECT 1.100000 1053.290000 1420.020000 1054.190000 ;
      RECT 0.000000 1047.480000 1420.020000 1053.290000 ;
      RECT 0.000000 1046.580000 1418.920000 1047.480000 ;
      RECT 0.000000 1045.040000 1420.020000 1046.580000 ;
      RECT 1.100000 1044.140000 1420.020000 1045.040000 ;
      RECT 0.000000 1038.330000 1420.020000 1044.140000 ;
      RECT 0.000000 1037.430000 1418.920000 1038.330000 ;
      RECT 0.000000 1035.890000 1420.020000 1037.430000 ;
      RECT 1.100000 1034.990000 1420.020000 1035.890000 ;
      RECT 0.000000 1029.180000 1420.020000 1034.990000 ;
      RECT 0.000000 1028.280000 1418.920000 1029.180000 ;
      RECT 0.000000 1027.350000 1420.020000 1028.280000 ;
      RECT 1.100000 1026.450000 1420.020000 1027.350000 ;
      RECT 0.000000 1020.030000 1420.020000 1026.450000 ;
      RECT 0.000000 1019.130000 1418.920000 1020.030000 ;
      RECT 0.000000 1018.200000 1420.020000 1019.130000 ;
      RECT 1.100000 1017.300000 1420.020000 1018.200000 ;
      RECT 0.000000 1011.490000 1420.020000 1017.300000 ;
      RECT 0.000000 1010.590000 1418.920000 1011.490000 ;
      RECT 0.000000 1009.660000 1420.020000 1010.590000 ;
      RECT 1.100000 1008.760000 1420.020000 1009.660000 ;
      RECT 0.000000 1002.340000 1420.020000 1008.760000 ;
      RECT 0.000000 1001.440000 1418.920000 1002.340000 ;
      RECT 0.000000 1000.510000 1420.020000 1001.440000 ;
      RECT 1.100000 999.610000 1420.020000 1000.510000 ;
      RECT 0.000000 993.190000 1420.020000 999.610000 ;
      RECT 0.000000 992.290000 1418.920000 993.190000 ;
      RECT 0.000000 991.360000 1420.020000 992.290000 ;
      RECT 1.100000 990.460000 1420.020000 991.360000 ;
      RECT 0.000000 984.040000 1420.020000 990.460000 ;
      RECT 0.000000 983.140000 1418.920000 984.040000 ;
      RECT 0.000000 982.820000 1420.020000 983.140000 ;
      RECT 1.100000 981.920000 1420.020000 982.820000 ;
      RECT 0.000000 974.890000 1420.020000 981.920000 ;
      RECT 0.000000 973.990000 1418.920000 974.890000 ;
      RECT 0.000000 973.670000 1420.020000 973.990000 ;
      RECT 1.100000 972.770000 1420.020000 973.670000 ;
      RECT 0.000000 965.740000 1420.020000 972.770000 ;
      RECT 0.000000 964.840000 1418.920000 965.740000 ;
      RECT 0.000000 964.520000 1420.020000 964.840000 ;
      RECT 1.100000 963.620000 1420.020000 964.520000 ;
      RECT 0.000000 956.590000 1420.020000 963.620000 ;
      RECT 0.000000 955.980000 1418.920000 956.590000 ;
      RECT 1.100000 955.690000 1418.920000 955.980000 ;
      RECT 1.100000 955.080000 1420.020000 955.690000 ;
      RECT 0.000000 947.440000 1420.020000 955.080000 ;
      RECT 0.000000 946.830000 1418.920000 947.440000 ;
      RECT 1.100000 946.540000 1418.920000 946.830000 ;
      RECT 1.100000 945.930000 1420.020000 946.540000 ;
      RECT 0.000000 938.290000 1420.020000 945.930000 ;
      RECT 1.100000 937.390000 1418.920000 938.290000 ;
      RECT 0.000000 929.140000 1420.020000 937.390000 ;
      RECT 1.100000 928.240000 1418.920000 929.140000 ;
      RECT 0.000000 919.990000 1420.020000 928.240000 ;
      RECT 1.100000 919.090000 1418.920000 919.990000 ;
      RECT 0.000000 911.450000 1420.020000 919.090000 ;
      RECT 1.100000 910.550000 1418.920000 911.450000 ;
      RECT 0.000000 902.300000 1420.020000 910.550000 ;
      RECT 1.100000 901.400000 1418.920000 902.300000 ;
      RECT 0.000000 893.150000 1420.020000 901.400000 ;
      RECT 1.100000 892.250000 1418.920000 893.150000 ;
      RECT 0.000000 884.610000 1420.020000 892.250000 ;
      RECT 1.100000 884.000000 1420.020000 884.610000 ;
      RECT 1.100000 883.710000 1418.920000 884.000000 ;
      RECT 0.000000 883.100000 1418.920000 883.710000 ;
      RECT 0.000000 875.460000 1420.020000 883.100000 ;
      RECT 1.100000 874.850000 1420.020000 875.460000 ;
      RECT 1.100000 874.560000 1418.920000 874.850000 ;
      RECT 0.000000 873.950000 1418.920000 874.560000 ;
      RECT 0.000000 866.920000 1420.020000 873.950000 ;
      RECT 1.100000 866.020000 1420.020000 866.920000 ;
      RECT 0.000000 865.700000 1420.020000 866.020000 ;
      RECT 0.000000 864.800000 1418.920000 865.700000 ;
      RECT 0.000000 857.770000 1420.020000 864.800000 ;
      RECT 1.100000 856.870000 1420.020000 857.770000 ;
      RECT 0.000000 856.550000 1420.020000 856.870000 ;
      RECT 0.000000 855.650000 1418.920000 856.550000 ;
      RECT 0.000000 848.620000 1420.020000 855.650000 ;
      RECT 1.100000 847.720000 1420.020000 848.620000 ;
      RECT 0.000000 847.400000 1420.020000 847.720000 ;
      RECT 0.000000 846.500000 1418.920000 847.400000 ;
      RECT 0.000000 840.080000 1420.020000 846.500000 ;
      RECT 1.100000 839.180000 1420.020000 840.080000 ;
      RECT 0.000000 838.250000 1420.020000 839.180000 ;
      RECT 0.000000 837.350000 1418.920000 838.250000 ;
      RECT 0.000000 830.930000 1420.020000 837.350000 ;
      RECT 1.100000 830.030000 1420.020000 830.930000 ;
      RECT 0.000000 829.100000 1420.020000 830.030000 ;
      RECT 0.000000 828.200000 1418.920000 829.100000 ;
      RECT 0.000000 821.780000 1420.020000 828.200000 ;
      RECT 1.100000 820.880000 1420.020000 821.780000 ;
      RECT 0.000000 819.950000 1420.020000 820.880000 ;
      RECT 0.000000 819.050000 1418.920000 819.950000 ;
      RECT 0.000000 813.240000 1420.020000 819.050000 ;
      RECT 1.100000 812.340000 1420.020000 813.240000 ;
      RECT 0.000000 811.410000 1420.020000 812.340000 ;
      RECT 0.000000 810.510000 1418.920000 811.410000 ;
      RECT 0.000000 804.090000 1420.020000 810.510000 ;
      RECT 1.100000 803.190000 1420.020000 804.090000 ;
      RECT 0.000000 802.260000 1420.020000 803.190000 ;
      RECT 0.000000 801.360000 1418.920000 802.260000 ;
      RECT 0.000000 794.940000 1420.020000 801.360000 ;
      RECT 1.100000 794.040000 1420.020000 794.940000 ;
      RECT 0.000000 793.110000 1420.020000 794.040000 ;
      RECT 0.000000 792.210000 1418.920000 793.110000 ;
      RECT 0.000000 786.400000 1420.020000 792.210000 ;
      RECT 1.100000 785.500000 1420.020000 786.400000 ;
      RECT 0.000000 783.960000 1420.020000 785.500000 ;
      RECT 0.000000 783.060000 1418.920000 783.960000 ;
      RECT 0.000000 777.250000 1420.020000 783.060000 ;
      RECT 1.100000 776.350000 1420.020000 777.250000 ;
      RECT 0.000000 774.810000 1420.020000 776.350000 ;
      RECT 0.000000 773.910000 1418.920000 774.810000 ;
      RECT 0.000000 768.710000 1420.020000 773.910000 ;
      RECT 1.100000 767.810000 1420.020000 768.710000 ;
      RECT 0.000000 765.660000 1420.020000 767.810000 ;
      RECT 0.000000 764.760000 1418.920000 765.660000 ;
      RECT 0.000000 759.560000 1420.020000 764.760000 ;
      RECT 1.100000 758.660000 1420.020000 759.560000 ;
      RECT 0.000000 756.510000 1420.020000 758.660000 ;
      RECT 0.000000 755.610000 1418.920000 756.510000 ;
      RECT 0.000000 750.410000 1420.020000 755.610000 ;
      RECT 1.100000 749.510000 1420.020000 750.410000 ;
      RECT 0.000000 747.360000 1420.020000 749.510000 ;
      RECT 0.000000 746.460000 1418.920000 747.360000 ;
      RECT 0.000000 741.870000 1420.020000 746.460000 ;
      RECT 1.100000 740.970000 1420.020000 741.870000 ;
      RECT 0.000000 738.210000 1420.020000 740.970000 ;
      RECT 0.000000 737.310000 1418.920000 738.210000 ;
      RECT 0.000000 732.720000 1420.020000 737.310000 ;
      RECT 1.100000 731.820000 1420.020000 732.720000 ;
      RECT 0.000000 729.060000 1420.020000 731.820000 ;
      RECT 0.000000 728.160000 1418.920000 729.060000 ;
      RECT 0.000000 723.570000 1420.020000 728.160000 ;
      RECT 1.100000 722.670000 1420.020000 723.570000 ;
      RECT 0.000000 719.910000 1420.020000 722.670000 ;
      RECT 0.000000 719.010000 1418.920000 719.910000 ;
      RECT 0.000000 715.030000 1420.020000 719.010000 ;
      RECT 1.100000 714.130000 1420.020000 715.030000 ;
      RECT 0.000000 710.760000 1420.020000 714.130000 ;
      RECT 0.000000 709.860000 1418.920000 710.760000 ;
      RECT 0.000000 705.880000 1420.020000 709.860000 ;
      RECT 1.100000 704.980000 1420.020000 705.880000 ;
      RECT 0.000000 702.220000 1420.020000 704.980000 ;
      RECT 0.000000 701.320000 1418.920000 702.220000 ;
      RECT 0.000000 697.340000 1420.020000 701.320000 ;
      RECT 1.100000 696.440000 1420.020000 697.340000 ;
      RECT 0.000000 693.070000 1420.020000 696.440000 ;
      RECT 0.000000 692.170000 1418.920000 693.070000 ;
      RECT 0.000000 688.190000 1420.020000 692.170000 ;
      RECT 1.100000 687.290000 1420.020000 688.190000 ;
      RECT 0.000000 683.920000 1420.020000 687.290000 ;
      RECT 0.000000 683.020000 1418.920000 683.920000 ;
      RECT 0.000000 679.040000 1420.020000 683.020000 ;
      RECT 1.100000 678.140000 1420.020000 679.040000 ;
      RECT 0.000000 674.770000 1420.020000 678.140000 ;
      RECT 0.000000 673.870000 1418.920000 674.770000 ;
      RECT 0.000000 670.500000 1420.020000 673.870000 ;
      RECT 1.100000 669.600000 1420.020000 670.500000 ;
      RECT 0.000000 665.620000 1420.020000 669.600000 ;
      RECT 0.000000 664.720000 1418.920000 665.620000 ;
      RECT 0.000000 661.350000 1420.020000 664.720000 ;
      RECT 1.100000 660.450000 1420.020000 661.350000 ;
      RECT 0.000000 656.470000 1420.020000 660.450000 ;
      RECT 0.000000 655.570000 1418.920000 656.470000 ;
      RECT 0.000000 652.200000 1420.020000 655.570000 ;
      RECT 1.100000 651.300000 1420.020000 652.200000 ;
      RECT 0.000000 647.320000 1420.020000 651.300000 ;
      RECT 0.000000 646.420000 1418.920000 647.320000 ;
      RECT 0.000000 643.660000 1420.020000 646.420000 ;
      RECT 1.100000 642.760000 1420.020000 643.660000 ;
      RECT 0.000000 638.170000 1420.020000 642.760000 ;
      RECT 0.000000 637.270000 1418.920000 638.170000 ;
      RECT 0.000000 634.510000 1420.020000 637.270000 ;
      RECT 1.100000 633.610000 1420.020000 634.510000 ;
      RECT 0.000000 629.020000 1420.020000 633.610000 ;
      RECT 0.000000 628.120000 1418.920000 629.020000 ;
      RECT 0.000000 625.970000 1420.020000 628.120000 ;
      RECT 1.100000 625.070000 1420.020000 625.970000 ;
      RECT 0.000000 619.870000 1420.020000 625.070000 ;
      RECT 0.000000 618.970000 1418.920000 619.870000 ;
      RECT 0.000000 616.820000 1420.020000 618.970000 ;
      RECT 1.100000 615.920000 1420.020000 616.820000 ;
      RECT 0.000000 610.720000 1420.020000 615.920000 ;
      RECT 0.000000 609.820000 1418.920000 610.720000 ;
      RECT 0.000000 607.670000 1420.020000 609.820000 ;
      RECT 1.100000 606.770000 1420.020000 607.670000 ;
      RECT 0.000000 602.180000 1420.020000 606.770000 ;
      RECT 0.000000 601.280000 1418.920000 602.180000 ;
      RECT 0.000000 599.130000 1420.020000 601.280000 ;
      RECT 1.100000 598.230000 1420.020000 599.130000 ;
      RECT 0.000000 593.030000 1420.020000 598.230000 ;
      RECT 0.000000 592.130000 1418.920000 593.030000 ;
      RECT 0.000000 589.980000 1420.020000 592.130000 ;
      RECT 1.100000 589.080000 1420.020000 589.980000 ;
      RECT 0.000000 583.880000 1420.020000 589.080000 ;
      RECT 0.000000 582.980000 1418.920000 583.880000 ;
      RECT 0.000000 580.830000 1420.020000 582.980000 ;
      RECT 1.100000 579.930000 1420.020000 580.830000 ;
      RECT 0.000000 574.730000 1420.020000 579.930000 ;
      RECT 0.000000 573.830000 1418.920000 574.730000 ;
      RECT 0.000000 572.290000 1420.020000 573.830000 ;
      RECT 1.100000 571.390000 1420.020000 572.290000 ;
      RECT 0.000000 565.580000 1420.020000 571.390000 ;
      RECT 0.000000 564.680000 1418.920000 565.580000 ;
      RECT 0.000000 563.140000 1420.020000 564.680000 ;
      RECT 1.100000 562.240000 1420.020000 563.140000 ;
      RECT 0.000000 556.430000 1420.020000 562.240000 ;
      RECT 0.000000 555.530000 1418.920000 556.430000 ;
      RECT 0.000000 553.990000 1420.020000 555.530000 ;
      RECT 1.100000 553.090000 1420.020000 553.990000 ;
      RECT 0.000000 547.280000 1420.020000 553.090000 ;
      RECT 0.000000 546.380000 1418.920000 547.280000 ;
      RECT 0.000000 545.450000 1420.020000 546.380000 ;
      RECT 1.100000 544.550000 1420.020000 545.450000 ;
      RECT 0.000000 538.130000 1420.020000 544.550000 ;
      RECT 0.000000 537.230000 1418.920000 538.130000 ;
      RECT 0.000000 536.300000 1420.020000 537.230000 ;
      RECT 1.100000 535.400000 1420.020000 536.300000 ;
      RECT 0.000000 528.980000 1420.020000 535.400000 ;
      RECT 0.000000 528.080000 1418.920000 528.980000 ;
      RECT 0.000000 527.760000 1420.020000 528.080000 ;
      RECT 1.100000 526.860000 1420.020000 527.760000 ;
      RECT 0.000000 519.830000 1420.020000 526.860000 ;
      RECT 0.000000 518.930000 1418.920000 519.830000 ;
      RECT 0.000000 518.610000 1420.020000 518.930000 ;
      RECT 1.100000 517.710000 1420.020000 518.610000 ;
      RECT 0.000000 510.680000 1420.020000 517.710000 ;
      RECT 0.000000 509.780000 1418.920000 510.680000 ;
      RECT 0.000000 509.460000 1420.020000 509.780000 ;
      RECT 1.100000 508.560000 1420.020000 509.460000 ;
      RECT 0.000000 502.140000 1420.020000 508.560000 ;
      RECT 0.000000 501.240000 1418.920000 502.140000 ;
      RECT 0.000000 500.920000 1420.020000 501.240000 ;
      RECT 1.100000 500.020000 1420.020000 500.920000 ;
      RECT 0.000000 492.990000 1420.020000 500.020000 ;
      RECT 0.000000 492.090000 1418.920000 492.990000 ;
      RECT 0.000000 491.770000 1420.020000 492.090000 ;
      RECT 1.100000 490.870000 1420.020000 491.770000 ;
      RECT 0.000000 483.840000 1420.020000 490.870000 ;
      RECT 0.000000 482.940000 1418.920000 483.840000 ;
      RECT 0.000000 482.620000 1420.020000 482.940000 ;
      RECT 1.100000 481.720000 1420.020000 482.620000 ;
      RECT 0.000000 474.690000 1420.020000 481.720000 ;
      RECT 0.000000 474.080000 1418.920000 474.690000 ;
      RECT 1.100000 473.790000 1418.920000 474.080000 ;
      RECT 1.100000 473.180000 1420.020000 473.790000 ;
      RECT 0.000000 465.540000 1420.020000 473.180000 ;
      RECT 0.000000 464.930000 1418.920000 465.540000 ;
      RECT 1.100000 464.640000 1418.920000 464.930000 ;
      RECT 1.100000 464.030000 1420.020000 464.640000 ;
      RECT 0.000000 456.390000 1420.020000 464.030000 ;
      RECT 1.100000 455.490000 1418.920000 456.390000 ;
      RECT 0.000000 447.240000 1420.020000 455.490000 ;
      RECT 1.100000 446.340000 1418.920000 447.240000 ;
      RECT 0.000000 438.090000 1420.020000 446.340000 ;
      RECT 1.100000 437.190000 1418.920000 438.090000 ;
      RECT 0.000000 429.550000 1420.020000 437.190000 ;
      RECT 1.100000 428.940000 1420.020000 429.550000 ;
      RECT 1.100000 428.650000 1418.920000 428.940000 ;
      RECT 0.000000 428.040000 1418.920000 428.650000 ;
      RECT 0.000000 420.400000 1420.020000 428.040000 ;
      RECT 1.100000 419.790000 1420.020000 420.400000 ;
      RECT 1.100000 419.500000 1418.920000 419.790000 ;
      RECT 0.000000 418.890000 1418.920000 419.500000 ;
      RECT 0.000000 411.250000 1420.020000 418.890000 ;
      RECT 1.100000 410.640000 1420.020000 411.250000 ;
      RECT 1.100000 410.350000 1418.920000 410.640000 ;
      RECT 0.000000 409.740000 1418.920000 410.350000 ;
      RECT 0.000000 402.710000 1420.020000 409.740000 ;
      RECT 1.100000 402.100000 1420.020000 402.710000 ;
      RECT 1.100000 401.810000 1418.920000 402.100000 ;
      RECT 0.000000 401.200000 1418.920000 401.810000 ;
      RECT 0.000000 393.560000 1420.020000 401.200000 ;
      RECT 1.100000 392.950000 1420.020000 393.560000 ;
      RECT 1.100000 392.660000 1418.920000 392.950000 ;
      RECT 0.000000 392.050000 1418.920000 392.660000 ;
      RECT 0.000000 385.020000 1420.020000 392.050000 ;
      RECT 1.100000 384.120000 1420.020000 385.020000 ;
      RECT 0.000000 383.800000 1420.020000 384.120000 ;
      RECT 0.000000 382.900000 1418.920000 383.800000 ;
      RECT 0.000000 375.870000 1420.020000 382.900000 ;
      RECT 1.100000 374.970000 1420.020000 375.870000 ;
      RECT 0.000000 374.650000 1420.020000 374.970000 ;
      RECT 0.000000 373.750000 1418.920000 374.650000 ;
      RECT 0.000000 366.720000 1420.020000 373.750000 ;
      RECT 1.100000 365.820000 1420.020000 366.720000 ;
      RECT 0.000000 365.500000 1420.020000 365.820000 ;
      RECT 0.000000 364.600000 1418.920000 365.500000 ;
      RECT 0.000000 358.180000 1420.020000 364.600000 ;
      RECT 1.100000 357.280000 1420.020000 358.180000 ;
      RECT 0.000000 356.350000 1420.020000 357.280000 ;
      RECT 0.000000 355.450000 1418.920000 356.350000 ;
      RECT 0.000000 349.030000 1420.020000 355.450000 ;
      RECT 1.100000 348.130000 1420.020000 349.030000 ;
      RECT 0.000000 347.200000 1420.020000 348.130000 ;
      RECT 0.000000 346.300000 1418.920000 347.200000 ;
      RECT 0.000000 339.880000 1420.020000 346.300000 ;
      RECT 1.100000 338.980000 1420.020000 339.880000 ;
      RECT 0.000000 338.050000 1420.020000 338.980000 ;
      RECT 0.000000 337.150000 1418.920000 338.050000 ;
      RECT 0.000000 331.340000 1420.020000 337.150000 ;
      RECT 1.100000 330.440000 1420.020000 331.340000 ;
      RECT 0.000000 328.900000 1420.020000 330.440000 ;
      RECT 0.000000 328.000000 1418.920000 328.900000 ;
      RECT 0.000000 322.190000 1420.020000 328.000000 ;
      RECT 1.100000 321.290000 1420.020000 322.190000 ;
      RECT 0.000000 319.750000 1420.020000 321.290000 ;
      RECT 0.000000 318.850000 1418.920000 319.750000 ;
      RECT 0.000000 313.650000 1420.020000 318.850000 ;
      RECT 1.100000 312.750000 1420.020000 313.650000 ;
      RECT 0.000000 310.600000 1420.020000 312.750000 ;
      RECT 0.000000 309.700000 1418.920000 310.600000 ;
      RECT 0.000000 304.500000 1420.020000 309.700000 ;
      RECT 1.100000 303.600000 1420.020000 304.500000 ;
      RECT 0.000000 302.060000 1420.020000 303.600000 ;
      RECT 0.000000 301.160000 1418.920000 302.060000 ;
      RECT 0.000000 295.350000 1420.020000 301.160000 ;
      RECT 1.100000 294.450000 1420.020000 295.350000 ;
      RECT 0.000000 292.910000 1420.020000 294.450000 ;
      RECT 0.000000 292.010000 1418.920000 292.910000 ;
      RECT 0.000000 286.810000 1420.020000 292.010000 ;
      RECT 1.100000 285.910000 1420.020000 286.810000 ;
      RECT 0.000000 283.760000 1420.020000 285.910000 ;
      RECT 0.000000 282.860000 1418.920000 283.760000 ;
      RECT 0.000000 277.660000 1420.020000 282.860000 ;
      RECT 1.100000 276.760000 1420.020000 277.660000 ;
      RECT 0.000000 274.610000 1420.020000 276.760000 ;
      RECT 0.000000 273.710000 1418.920000 274.610000 ;
      RECT 0.000000 268.510000 1420.020000 273.710000 ;
      RECT 1.100000 267.610000 1420.020000 268.510000 ;
      RECT 0.000000 265.460000 1420.020000 267.610000 ;
      RECT 0.000000 264.560000 1418.920000 265.460000 ;
      RECT 0.000000 259.970000 1420.020000 264.560000 ;
      RECT 1.100000 259.070000 1420.020000 259.970000 ;
      RECT 0.000000 256.310000 1420.020000 259.070000 ;
      RECT 0.000000 255.410000 1418.920000 256.310000 ;
      RECT 0.000000 250.820000 1420.020000 255.410000 ;
      RECT 1.100000 249.920000 1420.020000 250.820000 ;
      RECT 0.000000 247.160000 1420.020000 249.920000 ;
      RECT 0.000000 246.260000 1418.920000 247.160000 ;
      RECT 0.000000 241.670000 1420.020000 246.260000 ;
      RECT 1.100000 240.770000 1420.020000 241.670000 ;
      RECT 0.000000 238.010000 1420.020000 240.770000 ;
      RECT 0.000000 237.110000 1418.920000 238.010000 ;
      RECT 0.000000 233.130000 1420.020000 237.110000 ;
      RECT 1.100000 232.230000 1420.020000 233.130000 ;
      RECT 0.000000 228.860000 1420.020000 232.230000 ;
      RECT 0.000000 227.960000 1418.920000 228.860000 ;
      RECT 0.000000 223.980000 1420.020000 227.960000 ;
      RECT 1.100000 223.080000 1420.020000 223.980000 ;
      RECT 0.000000 219.710000 1420.020000 223.080000 ;
      RECT 0.000000 218.810000 1418.920000 219.710000 ;
      RECT 0.000000 215.440000 1420.020000 218.810000 ;
      RECT 1.100000 214.540000 1420.020000 215.440000 ;
      RECT 0.000000 210.560000 1420.020000 214.540000 ;
      RECT 0.000000 209.660000 1418.920000 210.560000 ;
      RECT 0.000000 206.290000 1420.020000 209.660000 ;
      RECT 1.100000 205.390000 1420.020000 206.290000 ;
      RECT 0.000000 202.020000 1420.020000 205.390000 ;
      RECT 0.000000 201.120000 1418.920000 202.020000 ;
      RECT 0.000000 197.140000 1420.020000 201.120000 ;
      RECT 1.100000 196.240000 1420.020000 197.140000 ;
      RECT 0.000000 192.870000 1420.020000 196.240000 ;
      RECT 0.000000 191.970000 1418.920000 192.870000 ;
      RECT 0.000000 188.600000 1420.020000 191.970000 ;
      RECT 1.100000 187.700000 1420.020000 188.600000 ;
      RECT 0.000000 183.720000 1420.020000 187.700000 ;
      RECT 0.000000 182.820000 1418.920000 183.720000 ;
      RECT 0.000000 179.450000 1420.020000 182.820000 ;
      RECT 1.100000 178.550000 1420.020000 179.450000 ;
      RECT 0.000000 174.570000 1420.020000 178.550000 ;
      RECT 0.000000 173.670000 1418.920000 174.570000 ;
      RECT 0.000000 170.300000 1420.020000 173.670000 ;
      RECT 1.100000 169.400000 1420.020000 170.300000 ;
      RECT 0.000000 165.420000 1420.020000 169.400000 ;
      RECT 0.000000 164.520000 1418.920000 165.420000 ;
      RECT 0.000000 161.760000 1420.020000 164.520000 ;
      RECT 1.100000 160.860000 1420.020000 161.760000 ;
      RECT 0.000000 156.270000 1420.020000 160.860000 ;
      RECT 0.000000 155.370000 1418.920000 156.270000 ;
      RECT 0.000000 152.610000 1420.020000 155.370000 ;
      RECT 1.100000 151.710000 1420.020000 152.610000 ;
      RECT 0.000000 147.120000 1420.020000 151.710000 ;
      RECT 0.000000 146.220000 1418.920000 147.120000 ;
      RECT 0.000000 144.070000 1420.020000 146.220000 ;
      RECT 1.100000 143.170000 1420.020000 144.070000 ;
      RECT 0.000000 137.970000 1420.020000 143.170000 ;
      RECT 0.000000 137.070000 1418.920000 137.970000 ;
      RECT 0.000000 134.920000 1420.020000 137.070000 ;
      RECT 1.100000 134.020000 1420.020000 134.920000 ;
      RECT 0.000000 128.820000 1420.020000 134.020000 ;
      RECT 0.000000 127.920000 1418.920000 128.820000 ;
      RECT 0.000000 125.770000 1420.020000 127.920000 ;
      RECT 1.100000 124.870000 1420.020000 125.770000 ;
      RECT 0.000000 119.670000 1420.020000 124.870000 ;
      RECT 0.000000 118.770000 1418.920000 119.670000 ;
      RECT 0.000000 117.230000 1420.020000 118.770000 ;
      RECT 1.100000 116.330000 1420.020000 117.230000 ;
      RECT 0.000000 110.520000 1420.020000 116.330000 ;
      RECT 0.000000 109.620000 1418.920000 110.520000 ;
      RECT 0.000000 108.080000 1420.020000 109.620000 ;
      RECT 1.100000 107.180000 1420.020000 108.080000 ;
      RECT 0.000000 101.980000 1420.020000 107.180000 ;
      RECT 0.000000 101.080000 1418.920000 101.980000 ;
      RECT 0.000000 98.930000 1420.020000 101.080000 ;
      RECT 1.100000 98.030000 1420.020000 98.930000 ;
      RECT 0.000000 92.830000 1420.020000 98.030000 ;
      RECT 0.000000 91.930000 1418.920000 92.830000 ;
      RECT 0.000000 90.390000 1420.020000 91.930000 ;
      RECT 1.100000 89.490000 1420.020000 90.390000 ;
      RECT 0.000000 83.680000 1420.020000 89.490000 ;
      RECT 0.000000 82.780000 1418.920000 83.680000 ;
      RECT 0.000000 81.240000 1420.020000 82.780000 ;
      RECT 1.100000 80.340000 1420.020000 81.240000 ;
      RECT 0.000000 74.530000 1420.020000 80.340000 ;
      RECT 0.000000 73.630000 1418.920000 74.530000 ;
      RECT 0.000000 72.700000 1420.020000 73.630000 ;
      RECT 1.100000 71.800000 1420.020000 72.700000 ;
      RECT 0.000000 65.380000 1420.020000 71.800000 ;
      RECT 0.000000 64.480000 1418.920000 65.380000 ;
      RECT 0.000000 63.550000 1420.020000 64.480000 ;
      RECT 1.100000 62.650000 1420.020000 63.550000 ;
      RECT 0.000000 56.230000 1420.020000 62.650000 ;
      RECT 0.000000 55.330000 1418.920000 56.230000 ;
      RECT 0.000000 54.400000 1420.020000 55.330000 ;
      RECT 1.100000 53.500000 1420.020000 54.400000 ;
      RECT 0.000000 47.080000 1420.020000 53.500000 ;
      RECT 0.000000 46.180000 1418.920000 47.080000 ;
      RECT 0.000000 45.860000 1420.020000 46.180000 ;
      RECT 1.100000 44.960000 1420.020000 45.860000 ;
      RECT 0.000000 37.930000 1420.020000 44.960000 ;
      RECT 0.000000 37.030000 1418.920000 37.930000 ;
      RECT 0.000000 36.710000 1420.020000 37.030000 ;
      RECT 1.100000 35.810000 1420.020000 36.710000 ;
      RECT 0.000000 28.780000 1420.020000 35.810000 ;
      RECT 0.000000 27.880000 1418.920000 28.780000 ;
      RECT 0.000000 27.560000 1420.020000 27.880000 ;
      RECT 1.100000 26.660000 1420.020000 27.560000 ;
      RECT 0.000000 19.630000 1420.020000 26.660000 ;
      RECT 0.000000 19.020000 1418.920000 19.630000 ;
      RECT 1.100000 18.730000 1418.920000 19.020000 ;
      RECT 1.100000 18.120000 1420.020000 18.730000 ;
      RECT 0.000000 10.480000 1420.020000 18.120000 ;
      RECT 0.000000 9.870000 1418.920000 10.480000 ;
      RECT 1.100000 9.580000 1418.920000 9.870000 ;
      RECT 1.100000 8.970000 1420.020000 9.580000 ;
      RECT 0.000000 8.360000 1420.020000 8.970000 ;
      RECT 1414.000000 5.760000 1420.020000 8.360000 ;
      RECT 0.000000 5.760000 6.020000 8.360000 ;
      RECT 0.000000 4.560000 1420.020000 5.760000 ;
      RECT 1417.800000 1.960000 1420.020000 4.560000 ;
      RECT 0.000000 1.960000 2.220000 4.560000 ;
      RECT 0.000000 1.940000 1420.020000 1.960000 ;
      RECT 1.100000 1.100000 1418.920000 1.940000 ;
      RECT 1411.500000 1.040000 1418.920000 1.100000 ;
      RECT 1.100000 1.040000 8.980000 1.100000 ;
      RECT 1411.500000 0.000000 1419.340000 1.040000 ;
      RECT 1402.760000 0.000000 1410.600000 1.100000 ;
      RECT 1393.560000 0.000000 1401.860000 1.100000 ;
      RECT 1384.820000 0.000000 1392.660000 1.100000 ;
      RECT 1375.620000 0.000000 1383.920000 1.100000 ;
      RECT 1366.880000 0.000000 1374.720000 1.100000 ;
      RECT 1358.140000 0.000000 1365.980000 1.100000 ;
      RECT 1348.940000 0.000000 1357.240000 1.100000 ;
      RECT 1340.200000 0.000000 1348.040000 1.100000 ;
      RECT 1331.000000 0.000000 1339.300000 1.100000 ;
      RECT 1322.260000 0.000000 1330.100000 1.100000 ;
      RECT 1313.520000 0.000000 1321.360000 1.100000 ;
      RECT 1304.320000 0.000000 1312.620000 1.100000 ;
      RECT 1295.580000 0.000000 1303.420000 1.100000 ;
      RECT 1286.380000 0.000000 1294.680000 1.100000 ;
      RECT 1277.640000 0.000000 1285.480000 1.100000 ;
      RECT 1268.900000 0.000000 1276.740000 1.100000 ;
      RECT 1259.700000 0.000000 1268.000000 1.100000 ;
      RECT 1250.960000 0.000000 1258.800000 1.100000 ;
      RECT 1241.760000 0.000000 1250.060000 1.100000 ;
      RECT 1233.020000 0.000000 1240.860000 1.100000 ;
      RECT 1224.280000 0.000000 1232.120000 1.100000 ;
      RECT 1215.080000 0.000000 1223.380000 1.100000 ;
      RECT 1206.340000 0.000000 1214.180000 1.100000 ;
      RECT 1197.140000 0.000000 1205.440000 1.100000 ;
      RECT 1188.400000 0.000000 1196.240000 1.100000 ;
      RECT 1179.200000 0.000000 1187.500000 1.100000 ;
      RECT 1170.460000 0.000000 1178.300000 1.100000 ;
      RECT 1161.720000 0.000000 1169.560000 1.100000 ;
      RECT 1152.520000 0.000000 1160.820000 1.100000 ;
      RECT 1143.780000 0.000000 1151.620000 1.100000 ;
      RECT 1134.580000 0.000000 1142.880000 1.100000 ;
      RECT 1125.840000 0.000000 1133.680000 1.100000 ;
      RECT 1117.100000 0.000000 1124.940000 1.100000 ;
      RECT 1107.900000 0.000000 1116.200000 1.100000 ;
      RECT 1099.160000 0.000000 1107.000000 1.100000 ;
      RECT 1089.960000 0.000000 1098.260000 1.100000 ;
      RECT 1081.220000 0.000000 1089.060000 1.100000 ;
      RECT 1072.480000 0.000000 1080.320000 1.100000 ;
      RECT 1063.280000 0.000000 1071.580000 1.100000 ;
      RECT 1054.540000 0.000000 1062.380000 1.100000 ;
      RECT 1045.340000 0.000000 1053.640000 1.100000 ;
      RECT 1036.600000 0.000000 1044.440000 1.100000 ;
      RECT 1027.860000 0.000000 1035.700000 1.100000 ;
      RECT 1018.660000 0.000000 1026.960000 1.100000 ;
      RECT 1009.920000 0.000000 1017.760000 1.100000 ;
      RECT 1000.720000 0.000000 1009.020000 1.100000 ;
      RECT 991.980000 0.000000 999.820000 1.100000 ;
      RECT 982.780000 0.000000 991.080000 1.100000 ;
      RECT 974.040000 0.000000 981.880000 1.100000 ;
      RECT 965.300000 0.000000 973.140000 1.100000 ;
      RECT 956.100000 0.000000 964.400000 1.100000 ;
      RECT 947.360000 0.000000 955.200000 1.100000 ;
      RECT 938.160000 0.000000 946.460000 1.100000 ;
      RECT 929.420000 0.000000 937.260000 1.100000 ;
      RECT 920.680000 0.000000 928.520000 1.100000 ;
      RECT 911.480000 0.000000 919.780000 1.100000 ;
      RECT 902.740000 0.000000 910.580000 1.100000 ;
      RECT 893.540000 0.000000 901.840000 1.100000 ;
      RECT 884.800000 0.000000 892.640000 1.100000 ;
      RECT 876.060000 0.000000 883.900000 1.100000 ;
      RECT 866.860000 0.000000 875.160000 1.100000 ;
      RECT 858.120000 0.000000 865.960000 1.100000 ;
      RECT 848.920000 0.000000 857.220000 1.100000 ;
      RECT 840.180000 0.000000 848.020000 1.100000 ;
      RECT 831.440000 0.000000 839.280000 1.100000 ;
      RECT 822.240000 0.000000 830.540000 1.100000 ;
      RECT 813.500000 0.000000 821.340000 1.100000 ;
      RECT 804.300000 0.000000 812.600000 1.100000 ;
      RECT 795.560000 0.000000 803.400000 1.100000 ;
      RECT 786.360000 0.000000 794.660000 1.100000 ;
      RECT 777.620000 0.000000 785.460000 1.100000 ;
      RECT 768.880000 0.000000 776.720000 1.100000 ;
      RECT 759.680000 0.000000 767.980000 1.100000 ;
      RECT 750.940000 0.000000 758.780000 1.100000 ;
      RECT 741.740000 0.000000 750.040000 1.100000 ;
      RECT 733.000000 0.000000 740.840000 1.100000 ;
      RECT 724.260000 0.000000 732.100000 1.100000 ;
      RECT 715.060000 0.000000 723.360000 1.100000 ;
      RECT 706.320000 0.000000 714.160000 1.100000 ;
      RECT 697.120000 0.000000 705.420000 1.100000 ;
      RECT 688.380000 0.000000 696.220000 1.100000 ;
      RECT 679.640000 0.000000 687.480000 1.100000 ;
      RECT 670.440000 0.000000 678.740000 1.100000 ;
      RECT 661.700000 0.000000 669.540000 1.100000 ;
      RECT 652.500000 0.000000 660.800000 1.100000 ;
      RECT 643.760000 0.000000 651.600000 1.100000 ;
      RECT 635.020000 0.000000 642.860000 1.100000 ;
      RECT 625.820000 0.000000 634.120000 1.100000 ;
      RECT 617.080000 0.000000 624.920000 1.100000 ;
      RECT 607.880000 0.000000 616.180000 1.100000 ;
      RECT 599.140000 0.000000 606.980000 1.100000 ;
      RECT 589.940000 0.000000 598.240000 1.100000 ;
      RECT 581.200000 0.000000 589.040000 1.100000 ;
      RECT 572.460000 0.000000 580.300000 1.100000 ;
      RECT 563.260000 0.000000 571.560000 1.100000 ;
      RECT 554.520000 0.000000 562.360000 1.100000 ;
      RECT 545.320000 0.000000 553.620000 1.100000 ;
      RECT 536.580000 0.000000 544.420000 1.100000 ;
      RECT 527.840000 0.000000 535.680000 1.100000 ;
      RECT 518.640000 0.000000 526.940000 1.100000 ;
      RECT 509.900000 0.000000 517.740000 1.100000 ;
      RECT 500.700000 0.000000 509.000000 1.100000 ;
      RECT 491.960000 0.000000 499.800000 1.100000 ;
      RECT 483.220000 0.000000 491.060000 1.100000 ;
      RECT 474.020000 0.000000 482.320000 1.100000 ;
      RECT 465.280000 0.000000 473.120000 1.100000 ;
      RECT 456.080000 0.000000 464.380000 1.100000 ;
      RECT 447.340000 0.000000 455.180000 1.100000 ;
      RECT 438.600000 0.000000 446.440000 1.100000 ;
      RECT 429.400000 0.000000 437.700000 1.100000 ;
      RECT 420.660000 0.000000 428.500000 1.100000 ;
      RECT 411.460000 0.000000 419.760000 1.100000 ;
      RECT 402.720000 0.000000 410.560000 1.100000 ;
      RECT 393.520000 0.000000 401.820000 1.100000 ;
      RECT 384.780000 0.000000 392.620000 1.100000 ;
      RECT 376.040000 0.000000 383.880000 1.100000 ;
      RECT 366.840000 0.000000 375.140000 1.100000 ;
      RECT 358.100000 0.000000 365.940000 1.100000 ;
      RECT 348.900000 0.000000 357.200000 1.100000 ;
      RECT 340.160000 0.000000 348.000000 1.100000 ;
      RECT 331.420000 0.000000 339.260000 1.100000 ;
      RECT 322.220000 0.000000 330.520000 1.100000 ;
      RECT 313.480000 0.000000 321.320000 1.100000 ;
      RECT 304.280000 0.000000 312.580000 1.100000 ;
      RECT 295.540000 0.000000 303.380000 1.100000 ;
      RECT 286.800000 0.000000 294.640000 1.100000 ;
      RECT 277.600000 0.000000 285.900000 1.100000 ;
      RECT 268.860000 0.000000 276.700000 1.100000 ;
      RECT 259.660000 0.000000 267.960000 1.100000 ;
      RECT 250.920000 0.000000 258.760000 1.100000 ;
      RECT 242.180000 0.000000 250.020000 1.100000 ;
      RECT 232.980000 0.000000 241.280000 1.100000 ;
      RECT 224.240000 0.000000 232.080000 1.100000 ;
      RECT 215.040000 0.000000 223.340000 1.100000 ;
      RECT 206.300000 0.000000 214.140000 1.100000 ;
      RECT 197.100000 0.000000 205.400000 1.100000 ;
      RECT 188.360000 0.000000 196.200000 1.100000 ;
      RECT 179.620000 0.000000 187.460000 1.100000 ;
      RECT 170.420000 0.000000 178.720000 1.100000 ;
      RECT 161.680000 0.000000 169.520000 1.100000 ;
      RECT 152.480000 0.000000 160.780000 1.100000 ;
      RECT 143.740000 0.000000 151.580000 1.100000 ;
      RECT 135.000000 0.000000 142.840000 1.100000 ;
      RECT 125.800000 0.000000 134.100000 1.100000 ;
      RECT 117.060000 0.000000 124.900000 1.100000 ;
      RECT 107.860000 0.000000 116.160000 1.100000 ;
      RECT 99.120000 0.000000 106.960000 1.100000 ;
      RECT 90.380000 0.000000 98.220000 1.100000 ;
      RECT 81.180000 0.000000 89.480000 1.100000 ;
      RECT 72.440000 0.000000 80.280000 1.100000 ;
      RECT 63.240000 0.000000 71.540000 1.100000 ;
      RECT 54.500000 0.000000 62.340000 1.100000 ;
      RECT 45.760000 0.000000 53.600000 1.100000 ;
      RECT 36.560000 0.000000 44.860000 1.100000 ;
      RECT 27.820000 0.000000 35.660000 1.100000 ;
      RECT 18.620000 0.000000 26.920000 1.100000 ;
      RECT 9.880000 0.000000 17.720000 1.100000 ;
      RECT 0.680000 0.000000 8.980000 1.040000 ;
    LAYER met4 ;
      RECT 0.000000 1415.840000 1420.020000 1419.840000 ;
      RECT 4.820000 1412.040000 1415.200000 1415.840000 ;
      RECT 1414.000000 5.760000 1415.200000 1412.040000 ;
      RECT 8.620000 5.760000 1411.400000 1412.040000 ;
      RECT 4.820000 5.760000 6.020000 1412.040000 ;
      RECT 1417.800000 1.960000 1420.020000 1415.840000 ;
      RECT 4.820000 1.960000 1415.200000 5.760000 ;
      RECT 0.000000 1.960000 2.220000 1415.840000 ;
      RECT 0.000000 0.000000 1420.020000 1.960000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 1420.020000 1419.840000 ;
  END
END soc_now_caravel_top

END LIBRARY
