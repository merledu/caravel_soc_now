magic
tech sky130A
magscale 1 2
timestamp 1669399178
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 397454 700476 397460 700528
rect 397512 700516 397518 700528
rect 459646 700516 459652 700528
rect 397512 700488 459652 700516
rect 397512 700476 397518 700488
rect 459646 700476 459652 700488
rect 459704 700476 459710 700528
rect 137830 700408 137836 700460
rect 137888 700448 137894 700460
rect 157978 700448 157984 700460
rect 137888 700420 157984 700448
rect 137888 700408 137894 700420
rect 157978 700408 157984 700420
rect 158036 700408 158042 700460
rect 255314 700408 255320 700460
rect 255372 700448 255378 700460
rect 332502 700448 332508 700460
rect 255372 700420 332508 700448
rect 255372 700408 255378 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 407114 700408 407120 700460
rect 407172 700448 407178 700460
rect 543458 700448 543464 700460
rect 407172 700420 543464 700448
rect 407172 700408 407178 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 8110 700340 8116 700392
rect 8168 700380 8174 700392
rect 131758 700380 131764 700392
rect 8168 700352 131764 700380
rect 8168 700340 8174 700352
rect 131758 700340 131764 700352
rect 131816 700340 131822 700392
rect 154114 700340 154120 700392
rect 154172 700380 154178 700392
rect 256694 700380 256700 700392
rect 154172 700352 256700 700380
rect 154172 700340 154178 700352
rect 256694 700340 256700 700352
rect 256752 700340 256758 700392
rect 267642 700340 267648 700392
rect 267700 700380 267706 700392
rect 436094 700380 436100 700392
rect 267700 700352 436100 700380
rect 267700 700340 267706 700352
rect 436094 700340 436100 700352
rect 436152 700340 436158 700392
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 227070 700312 227076 700324
rect 89220 700284 227076 700312
rect 89220 700272 89226 700284
rect 227070 700272 227076 700284
rect 227128 700272 227134 700324
rect 233970 700272 233976 700324
rect 234028 700312 234034 700324
rect 527174 700312 527180 700324
rect 234028 700284 527180 700312
rect 234028 700272 234034 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 306374 699700 306380 699712
rect 300176 699672 306380 699700
rect 300176 699660 300182 699672
rect 306374 699660 306380 699672
rect 306432 699660 306438 699712
rect 461670 699660 461676 699712
rect 461728 699700 461734 699712
rect 462314 699700 462320 699712
rect 461728 699672 462320 699700
rect 461728 699660 461734 699672
rect 462314 699660 462320 699672
rect 462372 699660 462378 699712
rect 465718 696940 465724 696992
rect 465776 696980 465782 696992
rect 580166 696980 580172 696992
rect 465776 696952 580172 696980
rect 465776 696940 465782 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 340874 683176 340880 683188
rect 3476 683148 340880 683176
rect 3476 683136 3482 683148
rect 340874 683136 340880 683148
rect 340932 683136 340938 683188
rect 498838 683136 498844 683188
rect 498896 683176 498902 683188
rect 580166 683176 580172 683188
rect 498896 683148 580172 683176
rect 498896 683136 498902 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 298094 670760 298100 670812
rect 298152 670800 298158 670812
rect 580166 670800 580172 670812
rect 298152 670772 580172 670800
rect 298152 670760 298158 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 452654 670732 452660 670744
rect 3568 670704 452660 670732
rect 3568 670692 3574 670704
rect 452654 670692 452660 670704
rect 452712 670692 452718 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 79318 656928 79324 656940
rect 3476 656900 79324 656928
rect 3476 656888 3482 656900
rect 79318 656888 79324 656900
rect 79376 656888 79382 656940
rect 502978 643084 502984 643136
rect 503036 643124 503042 643136
rect 580166 643124 580172 643136
rect 503036 643096 580172 643124
rect 503036 643084 503042 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 237374 630640 237380 630692
rect 237432 630680 237438 630692
rect 580166 630680 580172 630692
rect 237432 630652 580172 630680
rect 237432 630640 237438 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 314654 618304 314660 618316
rect 3200 618276 314660 618304
rect 3200 618264 3206 618276
rect 314654 618264 314660 618276
rect 314712 618264 314718 618316
rect 293954 616836 293960 616888
rect 294012 616876 294018 616888
rect 580166 616876 580172 616888
rect 294012 616848 580172 616876
rect 294012 616836 294018 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 485038 590656 485044 590708
rect 485096 590696 485102 590708
rect 579798 590696 579804 590708
rect 485096 590668 579804 590696
rect 485096 590656 485102 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 21358 579680 21364 579692
rect 3384 579652 21364 579680
rect 3384 579640 3390 579652
rect 21358 579640 21364 579652
rect 21416 579640 21422 579692
rect 3418 577464 3424 577516
rect 3476 577504 3482 577516
rect 453114 577504 453120 577516
rect 3476 577476 453120 577504
rect 3476 577464 3482 577476
rect 453114 577464 453120 577476
rect 453172 577464 453178 577516
rect 305454 574744 305460 574796
rect 305512 574784 305518 574796
rect 429194 574784 429200 574796
rect 305512 574756 429200 574784
rect 305512 574744 305518 574756
rect 429194 574744 429200 574756
rect 429252 574744 429258 574796
rect 234246 571956 234252 572008
rect 234304 571996 234310 572008
rect 412634 571996 412640 572008
rect 234304 571968 412640 571996
rect 234304 571956 234310 571968
rect 412634 571956 412640 571968
rect 412692 571956 412698 572008
rect 282914 570664 282920 570716
rect 282972 570704 282978 570716
rect 453022 570704 453028 570716
rect 282972 570676 453028 570704
rect 282972 570664 282978 570676
rect 453022 570664 453028 570676
rect 453080 570664 453086 570716
rect 234154 570596 234160 570648
rect 234212 570636 234218 570648
rect 580350 570636 580356 570648
rect 234212 570608 580356 570636
rect 234212 570596 234218 570608
rect 580350 570596 580356 570608
rect 580408 570596 580414 570648
rect 169754 566448 169760 566500
rect 169812 566488 169818 566500
rect 453206 566488 453212 566500
rect 169812 566460 453212 566488
rect 169812 566448 169818 566460
rect 453206 566448 453212 566460
rect 453264 566448 453270 566500
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 345382 565876 345388 565888
rect 3476 565848 345388 565876
rect 3476 565836 3482 565848
rect 345382 565836 345388 565848
rect 345440 565836 345446 565888
rect 234338 563728 234344 563780
rect 234396 563768 234402 563780
rect 347774 563768 347780 563780
rect 234396 563740 347780 563768
rect 234396 563728 234402 563740
rect 347774 563728 347780 563740
rect 347832 563728 347838 563780
rect 233142 563660 233148 563712
rect 233200 563700 233206 563712
rect 364334 563700 364340 563712
rect 233200 563672 364340 563700
rect 233200 563660 233206 563672
rect 364334 563660 364340 563672
rect 364392 563660 364398 563712
rect 406562 563048 406568 563100
rect 406620 563088 406626 563100
rect 579798 563088 579804 563100
rect 406620 563060 579804 563088
rect 406620 563048 406626 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 224310 562504 224316 562556
rect 224368 562544 224374 562556
rect 371786 562544 371792 562556
rect 224368 562516 371792 562544
rect 224368 562504 224374 562516
rect 371786 562504 371792 562516
rect 371844 562504 371850 562556
rect 215294 562436 215300 562488
rect 215352 562476 215358 562488
rect 426526 562476 426532 562488
rect 215352 562448 426532 562476
rect 215352 562436 215358 562448
rect 426526 562436 426532 562448
rect 426584 562436 426590 562488
rect 234522 562368 234528 562420
rect 234580 562408 234586 562420
rect 494054 562408 494060 562420
rect 234580 562380 494060 562408
rect 234580 562368 234586 562380
rect 494054 562368 494060 562380
rect 494112 562368 494118 562420
rect 104894 562300 104900 562352
rect 104952 562340 104958 562352
rect 456978 562340 456984 562352
rect 104952 562312 456984 562340
rect 104952 562300 104958 562312
rect 456978 562300 456984 562312
rect 457036 562300 457042 562352
rect 220446 562232 220452 562284
rect 220504 562272 220510 562284
rect 441614 562272 441620 562284
rect 220504 562244 441620 562272
rect 220504 562232 220510 562244
rect 441614 562232 441620 562244
rect 441672 562232 441678 562284
rect 106274 562164 106280 562216
rect 106332 562204 106338 562216
rect 340230 562204 340236 562216
rect 106332 562176 340236 562204
rect 106332 562164 106338 562176
rect 340230 562164 340236 562176
rect 340288 562164 340294 562216
rect 238754 562096 238760 562148
rect 238812 562136 238818 562148
rect 500954 562136 500960 562148
rect 238812 562108 500960 562136
rect 238812 562096 238818 562108
rect 500954 562096 500960 562108
rect 501012 562096 501018 562148
rect 253290 562028 253296 562080
rect 253348 562068 253354 562080
rect 531406 562068 531412 562080
rect 253348 562040 531412 562068
rect 253348 562028 253354 562040
rect 531406 562028 531412 562040
rect 531464 562028 531470 562080
rect 260374 561960 260380 562012
rect 260432 562000 260438 562012
rect 540974 562000 540980 562012
rect 260432 561972 540980 562000
rect 260432 561960 260438 561972
rect 540974 561960 540980 561972
rect 541032 561960 541038 562012
rect 279050 561892 279056 561944
rect 279108 561932 279114 561944
rect 572806 561932 572812 561944
rect 279108 561904 572812 561932
rect 279108 561892 279114 561904
rect 572806 561892 572812 561904
rect 572864 561892 572870 561944
rect 225966 561824 225972 561876
rect 226024 561864 226030 561876
rect 270678 561864 270684 561876
rect 226024 561836 270684 561864
rect 226024 561824 226030 561836
rect 270678 561824 270684 561836
rect 270736 561824 270742 561876
rect 273254 561824 273260 561876
rect 273312 561864 273318 561876
rect 576118 561864 576124 561876
rect 273312 561836 576124 561864
rect 273312 561824 273318 561836
rect 576118 561824 576124 561836
rect 576176 561824 576182 561876
rect 6914 561756 6920 561808
rect 6972 561796 6978 561808
rect 324314 561796 324320 561808
rect 6972 561768 324320 561796
rect 6972 561756 6978 561768
rect 324314 561756 324320 561768
rect 324372 561756 324378 561808
rect 241698 561688 241704 561740
rect 241756 561728 241762 561740
rect 569954 561728 569960 561740
rect 241756 561700 569960 561728
rect 241756 561688 241762 561700
rect 569954 561688 569960 561700
rect 570012 561688 570018 561740
rect 222838 561008 222844 561060
rect 222896 561048 222902 561060
rect 350534 561048 350540 561060
rect 222896 561020 350540 561048
rect 222896 561008 222902 561020
rect 350534 561008 350540 561020
rect 350592 561008 350598 561060
rect 252002 560940 252008 560992
rect 252060 560980 252066 560992
rect 558914 560980 558920 560992
rect 252060 560952 558920 560980
rect 252060 560940 252066 560952
rect 558914 560940 558920 560952
rect 558972 560940 558978 560992
rect 200758 560872 200764 560924
rect 200816 560912 200822 560924
rect 316034 560912 316040 560924
rect 200816 560884 316040 560912
rect 200816 560872 200822 560884
rect 316034 560872 316040 560884
rect 316092 560872 316098 560924
rect 329282 560872 329288 560924
rect 329340 560912 329346 560924
rect 483014 560912 483020 560924
rect 329340 560884 483020 560912
rect 329340 560872 329346 560884
rect 483014 560872 483020 560884
rect 483072 560872 483078 560924
rect 309318 560804 309324 560856
rect 309376 560844 309382 560856
rect 465810 560844 465816 560856
rect 309376 560816 465816 560844
rect 309376 560804 309382 560816
rect 465810 560804 465816 560816
rect 465868 560804 465874 560856
rect 227346 560736 227352 560788
rect 227404 560776 227410 560788
rect 271966 560776 271972 560788
rect 227404 560748 271972 560776
rect 227404 560736 227410 560748
rect 271966 560736 271972 560748
rect 272024 560736 272030 560788
rect 293218 560736 293224 560788
rect 293276 560776 293282 560788
rect 464522 560776 464528 560788
rect 293276 560748 464528 560776
rect 293276 560736 293282 560748
rect 464522 560736 464528 560748
rect 464580 560736 464586 560788
rect 206278 560668 206284 560720
rect 206336 560708 206342 560720
rect 382734 560708 382740 560720
rect 206336 560680 382740 560708
rect 206336 560668 206342 560680
rect 382734 560668 382740 560680
rect 382792 560668 382798 560720
rect 220170 560600 220176 560652
rect 220228 560640 220234 560652
rect 268102 560640 268108 560652
rect 220228 560612 268108 560640
rect 220228 560600 220234 560612
rect 268102 560600 268108 560612
rect 268160 560600 268166 560652
rect 302878 560600 302884 560652
rect 302936 560640 302942 560652
rect 480254 560640 480260 560652
rect 302936 560612 480260 560640
rect 302936 560600 302942 560612
rect 480254 560600 480260 560612
rect 480312 560600 480318 560652
rect 199378 560532 199384 560584
rect 199436 560572 199442 560584
rect 280338 560572 280344 560584
rect 199436 560544 280344 560572
rect 199436 560532 199442 560544
rect 280338 560532 280344 560544
rect 280396 560532 280402 560584
rect 300302 560532 300308 560584
rect 300360 560572 300366 560584
rect 487154 560572 487160 560584
rect 300360 560544 487160 560572
rect 300360 560532 300366 560544
rect 487154 560532 487160 560544
rect 487212 560532 487218 560584
rect 334434 560464 334440 560516
rect 334492 560504 334498 560516
rect 538858 560504 538864 560516
rect 334492 560476 538864 560504
rect 334492 560464 334498 560476
rect 538858 560464 538864 560476
rect 538916 560464 538922 560516
rect 244274 560396 244280 560448
rect 244332 560436 244338 560448
rect 507118 560436 507124 560448
rect 244332 560408 507124 560436
rect 244332 560396 244338 560408
rect 507118 560396 507124 560408
rect 507176 560396 507182 560448
rect 249794 560328 249800 560380
rect 249852 560368 249858 560380
rect 527818 560368 527824 560380
rect 249852 560340 527824 560368
rect 249852 560328 249858 560340
rect 527818 560328 527824 560340
rect 527876 560328 527882 560380
rect 8938 560260 8944 560312
rect 8996 560300 9002 560312
rect 445202 560300 445208 560312
rect 8996 560272 445208 560300
rect 8996 560260 9002 560272
rect 445202 560260 445208 560272
rect 445260 560260 445266 560312
rect 360930 559920 360936 559972
rect 360988 559960 360994 559972
rect 446582 559960 446588 559972
rect 360988 559932 446588 559960
rect 360988 559920 360994 559932
rect 446582 559920 446588 559932
rect 446640 559920 446646 559972
rect 234890 559852 234896 559904
rect 234948 559892 234954 559904
rect 368014 559892 368020 559904
rect 234948 559864 368020 559892
rect 234948 559852 234954 559864
rect 368014 559852 368020 559864
rect 368072 559852 368078 559904
rect 388622 559852 388628 559904
rect 388680 559892 388686 559904
rect 451734 559892 451740 559904
rect 388680 559864 451740 559892
rect 388680 559852 388686 559864
rect 451734 559852 451740 559864
rect 451792 559852 451798 559904
rect 232406 559784 232412 559836
rect 232464 559824 232470 559836
rect 393406 559824 393412 559836
rect 232464 559796 393412 559824
rect 232464 559784 232470 559796
rect 393406 559784 393412 559796
rect 393464 559784 393470 559836
rect 234706 559716 234712 559768
rect 234764 559756 234770 559768
rect 424042 559756 424048 559768
rect 234764 559728 424048 559756
rect 234764 559716 234770 559728
rect 424042 559716 424048 559728
rect 424100 559716 424106 559768
rect 223482 559648 223488 559700
rect 223540 559688 223546 559700
rect 245654 559688 245660 559700
rect 223540 559660 245660 559688
rect 223540 559648 223546 559660
rect 245654 559648 245660 559660
rect 245712 559648 245718 559700
rect 261662 559648 261668 559700
rect 261720 559688 261726 559700
rect 301682 559688 301688 559700
rect 261720 559660 301688 559688
rect 261720 559648 261726 559660
rect 301682 559648 301688 559660
rect 301740 559648 301746 559700
rect 419442 559648 419448 559700
rect 419500 559688 419506 559700
rect 459922 559688 459928 559700
rect 419500 559660 459928 559688
rect 419500 559648 419506 559660
rect 459922 559648 459928 559660
rect 459980 559648 459986 559700
rect 228358 559580 228364 559632
rect 228416 559620 228422 559632
rect 289446 559620 289452 559632
rect 228416 559592 289452 559620
rect 228416 559580 228422 559592
rect 289446 559580 289452 559592
rect 289504 559580 289510 559632
rect 416682 559580 416688 559632
rect 416740 559620 416746 559632
rect 461394 559620 461400 559632
rect 416740 559592 461400 559620
rect 416740 559580 416746 559592
rect 461394 559580 461400 559592
rect 461452 559580 461458 559632
rect 226794 559512 226800 559564
rect 226852 559552 226858 559564
rect 288434 559552 288440 559564
rect 226852 559524 288440 559552
rect 226852 559512 226858 559524
rect 288434 559512 288440 559524
rect 288492 559512 288498 559564
rect 414382 559512 414388 559564
rect 414440 559552 414446 559564
rect 460934 559552 460940 559564
rect 414440 559524 460940 559552
rect 414440 559512 414446 559524
rect 460934 559512 460940 559524
rect 460992 559512 460998 559564
rect 217318 559444 217324 559496
rect 217376 559484 217382 559496
rect 263042 559484 263048 559496
rect 217376 559456 263048 559484
rect 217376 559444 217382 559456
rect 263042 559444 263048 559456
rect 263100 559444 263106 559496
rect 274726 559444 274732 559496
rect 274784 559484 274790 559496
rect 362954 559484 362960 559496
rect 274784 559456 362960 559484
rect 274784 559444 274790 559456
rect 362954 559444 362960 559456
rect 363012 559444 363018 559496
rect 412450 559444 412456 559496
rect 412508 559484 412514 559496
rect 459002 559484 459008 559496
rect 412508 559456 459008 559484
rect 412508 559444 412514 559456
rect 459002 559444 459008 559456
rect 459060 559444 459066 559496
rect 229922 559376 229928 559428
rect 229980 559416 229986 559428
rect 322934 559416 322940 559428
rect 229980 559388 322940 559416
rect 229980 559376 229986 559388
rect 322934 559376 322940 559388
rect 322992 559376 322998 559428
rect 420822 559376 420828 559428
rect 420880 559416 420886 559428
rect 457070 559416 457076 559428
rect 420880 559388 457076 559416
rect 420880 559376 420886 559388
rect 457070 559376 457076 559388
rect 457128 559376 457134 559428
rect 167638 559308 167644 559360
rect 167696 559348 167702 559360
rect 292022 559348 292028 559360
rect 167696 559320 292028 559348
rect 167696 559308 167702 559320
rect 292022 559308 292028 559320
rect 292080 559308 292086 559360
rect 402146 559308 402152 559360
rect 402204 559348 402210 559360
rect 456886 559348 456892 559360
rect 402204 559320 456892 559348
rect 402204 559308 402210 559320
rect 456886 559308 456892 559320
rect 456944 559308 456950 559360
rect 224218 559240 224224 559292
rect 224276 559280 224282 559292
rect 354674 559280 354680 559292
rect 224276 559252 354680 559280
rect 224276 559240 224282 559252
rect 354674 559240 354680 559252
rect 354732 559240 354738 559292
rect 438210 559240 438216 559292
rect 438268 559280 438274 559292
rect 465350 559280 465356 559292
rect 438268 559252 465356 559280
rect 438268 559240 438274 559252
rect 465350 559240 465356 559252
rect 465408 559240 465414 559292
rect 367002 559172 367008 559224
rect 367060 559212 367066 559224
rect 389266 559212 389272 559224
rect 367060 559184 389272 559212
rect 367060 559172 367066 559184
rect 389266 559172 389272 559184
rect 389324 559172 389330 559224
rect 403434 559172 403440 559224
rect 403492 559212 403498 559224
rect 458358 559212 458364 559224
rect 403492 559184 458364 559212
rect 403492 559172 403498 559184
rect 458358 559172 458364 559184
rect 458416 559172 458422 559224
rect 235810 559104 235816 559156
rect 235868 559144 235874 559156
rect 378962 559144 378968 559156
rect 235868 559116 378968 559144
rect 235868 559104 235874 559116
rect 378962 559104 378968 559116
rect 379020 559104 379026 559156
rect 392486 559104 392492 559156
rect 392544 559144 392550 559156
rect 451642 559144 451648 559156
rect 392544 559116 451648 559144
rect 392544 559104 392550 559116
rect 451642 559104 451648 559116
rect 451700 559104 451706 559156
rect 228450 559036 228456 559088
rect 228508 559076 228514 559088
rect 377674 559076 377680 559088
rect 228508 559048 377680 559076
rect 228508 559036 228514 559048
rect 377674 559036 377680 559048
rect 377732 559036 377738 559088
rect 378778 559036 378784 559088
rect 378836 559076 378842 559088
rect 430574 559076 430580 559088
rect 378836 559048 430580 559076
rect 378836 559036 378842 559048
rect 430574 559036 430580 559048
rect 430632 559036 430638 559088
rect 432414 559036 432420 559088
rect 432472 559076 432478 559088
rect 464062 559076 464068 559088
rect 432472 559048 464068 559076
rect 432472 559036 432478 559048
rect 464062 559036 464068 559048
rect 464120 559036 464126 559088
rect 235902 558968 235908 559020
rect 235960 559008 235966 559020
rect 261754 559008 261760 559020
rect 235960 558980 261760 559008
rect 235960 558968 235966 558980
rect 261754 558968 261760 558980
rect 261812 558968 261818 559020
rect 262858 558968 262864 559020
rect 262916 559008 262922 559020
rect 274634 559008 274640 559020
rect 262916 558980 274640 559008
rect 262916 558968 262922 558980
rect 274634 558968 274640 558980
rect 274692 558968 274698 559020
rect 398282 558968 398288 559020
rect 398340 559008 398346 559020
rect 462406 559008 462412 559020
rect 398340 558980 462412 559008
rect 398340 558968 398346 558980
rect 462406 558968 462412 558980
rect 462464 558968 462470 559020
rect 232774 558900 232780 558952
rect 232832 558940 232838 558952
rect 265618 558940 265624 558952
rect 232832 558912 265624 558940
rect 232832 558900 232838 558912
rect 265618 558900 265624 558912
rect 265676 558900 265682 558952
rect 393314 558900 393320 558952
rect 393372 558940 393378 558952
rect 421466 558940 421472 558952
rect 393372 558912 421472 558940
rect 393372 558900 393378 558912
rect 421466 558900 421472 558912
rect 421524 558900 421530 558952
rect 423398 558900 423404 558952
rect 423456 558940 423462 558952
rect 469858 558940 469864 558952
rect 423456 558912 469864 558940
rect 423456 558900 423462 558912
rect 469858 558900 469864 558912
rect 469916 558900 469922 558952
rect 225598 558424 225604 558476
rect 225656 558464 225662 558476
rect 284294 558464 284300 558476
rect 225656 558436 284300 558464
rect 225656 558424 225662 558436
rect 284294 558424 284300 558436
rect 284352 558424 284358 558476
rect 225414 558356 225420 558408
rect 225472 558396 225478 558408
rect 287054 558396 287060 558408
rect 225472 558368 287060 558396
rect 225472 558356 225478 558368
rect 287054 558356 287060 558368
rect 287112 558356 287118 558408
rect 155954 558288 155960 558340
rect 156012 558328 156018 558340
rect 274726 558328 274732 558340
rect 156012 558300 274732 558328
rect 156012 558288 156018 558300
rect 274726 558288 274732 558300
rect 274784 558288 274790 558340
rect 46934 558220 46940 558272
rect 46992 558260 46998 558272
rect 262858 558260 262864 558272
rect 46992 558232 262864 558260
rect 46992 558220 46998 558232
rect 262858 558220 262864 558232
rect 262916 558220 262922 558272
rect 343542 558220 343548 558272
rect 343600 558260 343606 558272
rect 453298 558260 453304 558272
rect 343600 558232 453304 558260
rect 343600 558220 343606 558232
rect 453298 558220 453304 558232
rect 453356 558220 453362 558272
rect 3418 558152 3424 558204
rect 3476 558192 3482 558204
rect 378778 558192 378784 558204
rect 3476 558164 378784 558192
rect 3476 558152 3482 558164
rect 378778 558152 378784 558164
rect 378836 558152 378842 558204
rect 400858 558152 400864 558204
rect 400916 558192 400922 558204
rect 481726 558192 481732 558204
rect 400916 558164 481732 558192
rect 400916 558152 400922 558164
rect 481726 558152 481732 558164
rect 481784 558152 481790 558204
rect 233878 558084 233884 558136
rect 233936 558124 233942 558136
rect 320358 558124 320364 558136
rect 233936 558096 320364 558124
rect 233936 558084 233942 558096
rect 320358 558084 320364 558096
rect 320416 558084 320422 558136
rect 349982 558084 349988 558136
rect 350040 558124 350046 558136
rect 460198 558124 460204 558136
rect 350040 558096 460204 558124
rect 350040 558084 350046 558096
rect 460198 558084 460204 558096
rect 460256 558084 460262 558136
rect 232866 558016 232872 558068
rect 232924 558056 232930 558068
rect 328086 558056 328092 558068
rect 232924 558028 328092 558056
rect 232924 558016 232930 558028
rect 328086 558016 328092 558028
rect 328144 558016 328150 558068
rect 449802 558016 449808 558068
rect 449860 558056 449866 558068
rect 472618 558056 472624 558068
rect 449860 558028 472624 558056
rect 449860 558016 449866 558028
rect 472618 558016 472624 558028
rect 472676 558016 472682 558068
rect 187694 557948 187700 558000
rect 187752 557988 187758 558000
rect 356422 557988 356428 558000
rect 187752 557960 356428 557988
rect 187752 557948 187758 557960
rect 356422 557948 356428 557960
rect 356480 557948 356486 558000
rect 404722 557948 404728 558000
rect 404780 557988 404786 558000
rect 503714 557988 503720 558000
rect 404780 557960 503720 557988
rect 404780 557948 404786 557960
rect 503714 557948 503720 557960
rect 503772 557948 503778 558000
rect 136634 557880 136640 557932
rect 136692 557920 136698 557932
rect 317782 557920 317788 557932
rect 136692 557892 317788 557920
rect 136692 557880 136698 557892
rect 317782 557880 317788 557892
rect 317840 557880 317846 557932
rect 344830 557880 344836 557932
rect 344888 557920 344894 557932
rect 466454 557920 466460 557932
rect 344888 557892 466460 557920
rect 344888 557880 344894 557892
rect 466454 557880 466460 557892
rect 466512 557880 466518 557932
rect 92474 557812 92480 557864
rect 92532 557852 92538 557864
rect 285674 557852 285680 557864
rect 92532 557824 285680 557852
rect 92532 557812 92538 557824
rect 285674 557812 285680 557824
rect 285732 557812 285738 557864
rect 391198 557812 391204 557864
rect 391256 557852 391262 557864
rect 524414 557852 524420 557864
rect 391256 557824 524420 557852
rect 391256 557812 391262 557824
rect 524414 557812 524420 557824
rect 524472 557812 524478 557864
rect 15194 557744 15200 557796
rect 15252 557784 15258 557796
rect 259454 557784 259460 557796
rect 15252 557756 259460 557784
rect 15252 557744 15258 557756
rect 259454 557744 259460 557756
rect 259512 557744 259518 557796
rect 308766 557744 308772 557796
rect 308824 557784 308830 557796
rect 465166 557784 465172 557796
rect 308824 557756 465172 557784
rect 308824 557744 308830 557756
rect 465166 557744 465172 557756
rect 465224 557744 465230 557796
rect 241146 557676 241152 557728
rect 241204 557716 241210 557728
rect 492674 557716 492680 557728
rect 241204 557688 492680 557716
rect 241204 557676 241210 557688
rect 492674 557676 492680 557688
rect 492732 557676 492738 557728
rect 162854 557608 162860 557660
rect 162912 557648 162918 557660
rect 433702 557648 433708 557660
rect 162912 557620 433708 557648
rect 162912 557608 162918 557620
rect 433702 557608 433708 557620
rect 433760 557608 433766 557660
rect 443362 557608 443368 557660
rect 443420 557648 443426 557660
rect 496814 557648 496820 557660
rect 443420 557620 496820 557648
rect 443420 557608 443426 557620
rect 496814 557608 496820 557620
rect 496872 557608 496878 557660
rect 126974 557540 126980 557592
rect 127032 557580 127038 557592
rect 405366 557580 405372 557592
rect 127032 557552 405372 557580
rect 127032 557540 127038 557552
rect 405366 557540 405372 557552
rect 405424 557540 405430 557592
rect 435634 557540 435640 557592
rect 435692 557580 435698 557592
rect 565814 557580 565820 557592
rect 435692 557552 565820 557580
rect 435692 557540 435698 557552
rect 565814 557540 565820 557552
rect 565872 557540 565878 557592
rect 197354 557132 197360 557184
rect 197412 557172 197418 557184
rect 353294 557172 353300 557184
rect 197412 557144 353300 557172
rect 197412 557132 197418 557144
rect 353294 557132 353300 557144
rect 353352 557132 353358 557184
rect 143534 557064 143540 557116
rect 143592 557104 143598 557116
rect 369302 557104 369308 557116
rect 143592 557076 369308 557104
rect 143592 557064 143598 557076
rect 369302 557064 369308 557076
rect 369360 557064 369366 557116
rect 386046 557064 386052 557116
rect 386104 557104 386110 557116
rect 453574 557104 453580 557116
rect 386104 557076 453580 557104
rect 386104 557064 386110 557076
rect 453574 557064 453580 557076
rect 453632 557064 453638 557116
rect 127066 556996 127072 557048
rect 127124 557036 127130 557048
rect 366726 557036 366732 557048
rect 127124 557008 366732 557036
rect 127124 556996 127130 557008
rect 366726 556996 366732 557008
rect 366784 556996 366790 557048
rect 376662 556996 376668 557048
rect 376720 557036 376726 557048
rect 451550 557036 451556 557048
rect 376720 557008 451556 557036
rect 376720 556996 376726 557008
rect 451550 556996 451556 557008
rect 451608 556996 451614 557048
rect 226150 556928 226156 556980
rect 226208 556968 226214 556980
rect 266906 556968 266912 556980
rect 226208 556940 266912 556968
rect 226208 556928 226214 556940
rect 266906 556928 266912 556940
rect 266964 556928 266970 556980
rect 387334 556928 387340 556980
rect 387392 556968 387398 556980
rect 469214 556968 469220 556980
rect 387392 556940 469220 556968
rect 387392 556928 387398 556940
rect 469214 556928 469220 556940
rect 469272 556928 469278 556980
rect 175274 556860 175280 556912
rect 175332 556900 175338 556912
rect 393314 556900 393320 556912
rect 175332 556872 393320 556900
rect 175332 556860 175338 556872
rect 393314 556860 393320 556872
rect 393372 556860 393378 556912
rect 425974 556860 425980 556912
rect 426032 556900 426038 556912
rect 495434 556900 495440 556912
rect 426032 556872 495440 556900
rect 426032 556860 426038 556872
rect 495434 556860 495440 556872
rect 495492 556860 495498 556912
rect 3510 556792 3516 556844
rect 3568 556832 3574 556844
rect 360930 556832 360936 556844
rect 3568 556804 360936 556832
rect 3568 556792 3574 556804
rect 360930 556792 360936 556804
rect 360988 556792 360994 556844
rect 370912 556792 370918 556844
rect 370970 556832 370976 556844
rect 462498 556832 462504 556844
rect 370970 556804 462504 556832
rect 370970 556792 370976 556804
rect 462498 556792 462504 556804
rect 462556 556792 462562 556844
rect 207014 556724 207020 556776
rect 207072 556764 207078 556776
rect 248552 556764 248558 556776
rect 207072 556736 248558 556764
rect 207072 556724 207078 556736
rect 248552 556724 248558 556736
rect 248610 556724 248616 556776
rect 333560 556724 333566 556776
rect 333618 556764 333624 556776
rect 461118 556764 461124 556776
rect 333618 556736 461124 556764
rect 333618 556724 333624 556736
rect 461118 556724 461124 556736
rect 461176 556724 461182 556776
rect 218054 556656 218060 556708
rect 218112 556696 218118 556708
rect 321646 556696 321652 556708
rect 218112 556668 321652 556696
rect 218112 556656 218118 556668
rect 321646 556656 321652 556668
rect 321704 556656 321710 556708
rect 332502 556656 332508 556708
rect 332560 556696 332566 556708
rect 462590 556696 462596 556708
rect 332560 556668 462596 556696
rect 332560 556656 332566 556668
rect 462590 556656 462596 556668
rect 462648 556656 462654 556708
rect 227622 556588 227628 556640
rect 227680 556628 227686 556640
rect 269482 556628 269488 556640
rect 227680 556600 269488 556628
rect 227680 556588 227686 556600
rect 269482 556588 269488 556600
rect 269540 556588 269546 556640
rect 312630 556588 312636 556640
rect 312688 556628 312694 556640
rect 459554 556628 459560 556640
rect 312688 556600 459560 556628
rect 312688 556588 312694 556600
rect 459554 556588 459560 556600
rect 459612 556588 459618 556640
rect 233786 556520 233792 556572
rect 233844 556560 233850 556572
rect 234890 556560 234896 556572
rect 233844 556532 234896 556560
rect 233844 556520 233850 556532
rect 234890 556520 234896 556532
rect 234948 556520 234954 556572
rect 339494 556520 339500 556572
rect 339552 556560 339558 556572
rect 453666 556560 453672 556572
rect 339552 556532 453672 556560
rect 339552 556520 339558 556532
rect 453666 556520 453672 556532
rect 453724 556520 453730 556572
rect 193306 556452 193312 556504
rect 193364 556492 193370 556504
rect 358998 556492 359004 556504
rect 193364 556464 359004 556492
rect 193364 556452 193370 556464
rect 358998 556452 359004 556464
rect 359056 556452 359062 556504
rect 360930 556452 360936 556504
rect 360988 556492 360994 556504
rect 518894 556492 518900 556504
rect 360988 556464 518900 556492
rect 360988 556452 360994 556464
rect 518894 556452 518900 556464
rect 518952 556452 518958 556504
rect 227714 556384 227720 556436
rect 227772 556424 227778 556436
rect 283006 556424 283012 556436
rect 227772 556396 283012 556424
rect 227772 556384 227778 556396
rect 283006 556384 283012 556396
rect 283064 556384 283070 556436
rect 291194 556384 291200 556436
rect 291252 556424 291258 556436
rect 461026 556424 461032 556436
rect 291252 556396 461032 556424
rect 291252 556384 291258 556396
rect 461026 556384 461032 556396
rect 461084 556384 461090 556436
rect 193214 556316 193220 556368
rect 193272 556356 193278 556368
rect 276014 556356 276020 556368
rect 193272 556328 276020 556356
rect 193272 556316 193278 556328
rect 276014 556316 276020 556328
rect 276072 556316 276078 556368
rect 296438 556316 296444 556368
rect 296496 556356 296502 556368
rect 511994 556356 512000 556368
rect 296496 556328 512000 556356
rect 296496 556316 296502 556328
rect 511994 556316 512000 556328
rect 512052 556316 512058 556368
rect 226978 556248 226984 556300
rect 227036 556288 227042 556300
rect 247034 556288 247040 556300
rect 227036 556260 247040 556288
rect 227036 556248 227042 556260
rect 247034 556248 247040 556260
rect 247092 556248 247098 556300
rect 395706 556248 395712 556300
rect 395764 556288 395770 556300
rect 513374 556288 513380 556300
rect 395764 556260 513380 556288
rect 395764 556248 395770 556260
rect 513374 556248 513380 556260
rect 513432 556248 513438 556300
rect 226058 556180 226064 556232
rect 226116 556220 226122 556232
rect 254670 556220 254676 556232
rect 226116 556192 254676 556220
rect 226116 556180 226122 556192
rect 254670 556180 254676 556192
rect 254728 556180 254734 556232
rect 399570 556180 399576 556232
rect 399628 556220 399634 556232
rect 571978 556220 571984 556232
rect 399628 556192 571984 556220
rect 399628 556180 399634 556192
rect 571978 556180 571984 556192
rect 572036 556180 572042 556232
rect 235810 556084 235816 556096
rect 219406 556056 235816 556084
rect 117314 555704 117320 555756
rect 117372 555744 117378 555756
rect 219406 555744 219434 556056
rect 235810 556044 235816 556056
rect 235868 556044 235874 556096
rect 235902 556044 235908 556096
rect 235960 556044 235966 556096
rect 261662 556084 261668 556096
rect 258046 556056 261668 556084
rect 234706 555976 234712 556028
rect 234764 556016 234770 556028
rect 235920 556016 235948 556044
rect 234764 555988 235948 556016
rect 234764 555976 234770 555988
rect 117372 555716 219434 555744
rect 117372 555704 117378 555716
rect 114554 555636 114560 555688
rect 114612 555676 114618 555688
rect 234798 555676 234804 555688
rect 114612 555648 234804 555676
rect 114612 555636 114618 555648
rect 234798 555636 234804 555648
rect 234856 555636 234862 555688
rect 107654 555568 107660 555620
rect 107712 555608 107718 555620
rect 234706 555608 234712 555620
rect 107712 555580 234712 555608
rect 107712 555568 107718 555580
rect 234706 555568 234712 555580
rect 234764 555568 234770 555620
rect 86954 555500 86960 555552
rect 87012 555540 87018 555552
rect 234890 555540 234896 555552
rect 87012 555512 234896 555540
rect 87012 555500 87018 555512
rect 234890 555500 234896 555512
rect 234948 555500 234954 555552
rect 3602 555432 3608 555484
rect 3660 555472 3666 555484
rect 258046 555472 258074 556056
rect 261662 556044 261668 556056
rect 261720 556044 261726 556096
rect 364794 556044 364800 556096
rect 364852 556084 364858 556096
rect 364852 556056 373994 556084
rect 364852 556044 364858 556056
rect 3660 555444 258074 555472
rect 3660 555432 3666 555444
rect 223298 554752 223304 554804
rect 223356 554792 223362 554804
rect 232038 554792 232044 554804
rect 223356 554764 232044 554792
rect 223356 554752 223362 554764
rect 232038 554752 232044 554764
rect 232096 554752 232102 554804
rect 373966 554792 373994 556056
rect 451642 555432 451648 555484
rect 451700 555472 451706 555484
rect 580350 555472 580356 555484
rect 451700 555444 580356 555472
rect 451700 555432 451706 555444
rect 580350 555432 580356 555444
rect 580408 555432 580414 555484
rect 454034 554792 454040 554804
rect 373966 554764 454040 554792
rect 454034 554752 454040 554764
rect 454092 554752 454098 554804
rect 211798 554072 211804 554124
rect 211856 554112 211862 554124
rect 233050 554112 233056 554124
rect 211856 554084 233056 554112
rect 211856 554072 211862 554084
rect 233050 554072 233056 554084
rect 233108 554072 233114 554124
rect 118694 554004 118700 554056
rect 118752 554044 118758 554056
rect 233786 554044 233792 554056
rect 118752 554016 233792 554044
rect 118752 554004 118758 554016
rect 233786 554004 233792 554016
rect 233844 554004 233850 554056
rect 451734 554004 451740 554056
rect 451792 554044 451798 554056
rect 580258 554044 580264 554056
rect 451792 554016 580264 554044
rect 451792 554004 451798 554016
rect 580258 554004 580264 554016
rect 580316 554004 580322 554056
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 10318 553432 10324 553444
rect 3384 553404 10324 553432
rect 3384 553392 3390 553404
rect 10318 553392 10324 553404
rect 10376 553392 10382 553444
rect 223390 553392 223396 553444
rect 223448 553432 223454 553444
rect 232038 553432 232044 553444
rect 223448 553404 232044 553432
rect 223448 553392 223454 553404
rect 232038 553392 232044 553404
rect 232096 553392 232102 553444
rect 453942 553392 453948 553444
rect 454000 553432 454006 553444
rect 468570 553432 468576 553444
rect 454000 553404 468576 553432
rect 454000 553392 454006 553404
rect 468570 553392 468576 553404
rect 468628 553392 468634 553444
rect 59998 552032 60004 552084
rect 60056 552072 60062 552084
rect 232038 552072 232044 552084
rect 60056 552044 232044 552072
rect 60056 552032 60062 552044
rect 232038 552032 232044 552044
rect 232096 552032 232102 552084
rect 452930 551284 452936 551336
rect 452988 551324 452994 551336
rect 574094 551324 574100 551336
rect 452988 551296 574100 551324
rect 452988 551284 452994 551296
rect 574094 551284 574100 551296
rect 574152 551284 574158 551336
rect 160094 550604 160100 550656
rect 160152 550644 160158 550656
rect 232038 550644 232044 550656
rect 160152 550616 232044 550644
rect 160152 550604 160158 550616
rect 232038 550604 232044 550616
rect 232096 550604 232102 550656
rect 2774 549856 2780 549908
rect 2832 549896 2838 549908
rect 232774 549896 232780 549908
rect 2832 549868 232780 549896
rect 2832 549856 2838 549868
rect 232774 549856 232780 549868
rect 232832 549856 232838 549908
rect 453390 549448 453396 549500
rect 453448 549488 453454 549500
rect 455690 549488 455696 549500
rect 453448 549460 455696 549488
rect 453448 549448 453454 549460
rect 455690 549448 455696 549460
rect 455748 549448 455754 549500
rect 104894 548496 104900 548548
rect 104952 548536 104958 548548
rect 232406 548536 232412 548548
rect 104952 548508 232412 548536
rect 104952 548496 104958 548508
rect 232406 548496 232412 548508
rect 232464 548496 232470 548548
rect 26234 547136 26240 547188
rect 26292 547176 26298 547188
rect 232774 547176 232780 547188
rect 26292 547148 232780 547176
rect 26292 547136 26298 547148
rect 232774 547136 232780 547148
rect 232832 547136 232838 547188
rect 453942 546524 453948 546576
rect 454000 546564 454006 546576
rect 457622 546564 457628 546576
rect 454000 546536 457628 546564
rect 454000 546524 454006 546536
rect 457622 546524 457628 546536
rect 457680 546524 457686 546576
rect 176654 545096 176660 545148
rect 176712 545136 176718 545148
rect 232038 545136 232044 545148
rect 176712 545108 232044 545136
rect 176712 545096 176718 545108
rect 232038 545096 232044 545108
rect 232096 545096 232102 545148
rect 453942 545096 453948 545148
rect 454000 545136 454006 545148
rect 536834 545136 536840 545148
rect 454000 545108 536840 545136
rect 454000 545096 454006 545108
rect 536834 545096 536840 545108
rect 536892 545096 536898 545148
rect 60734 544348 60740 544400
rect 60792 544388 60798 544400
rect 232590 544388 232596 544400
rect 60792 544360 232596 544388
rect 60792 544348 60798 544360
rect 232590 544348 232596 544360
rect 232648 544348 232654 544400
rect 453574 544008 453580 544060
rect 453632 544048 453638 544060
rect 455598 544048 455604 544060
rect 453632 544020 455604 544048
rect 453632 544008 453638 544020
rect 455598 544008 455604 544020
rect 455656 544008 455662 544060
rect 67634 542988 67640 543040
rect 67692 543028 67698 543040
rect 228450 543028 228456 543040
rect 67692 543000 228456 543028
rect 67692 542988 67698 543000
rect 228450 542988 228456 543000
rect 228508 542988 228514 543040
rect 453942 542376 453948 542428
rect 454000 542416 454006 542428
rect 468478 542416 468484 542428
rect 454000 542388 468484 542416
rect 454000 542376 454006 542388
rect 468478 542376 468484 542388
rect 468536 542376 468542 542428
rect 233050 541220 233056 541272
rect 233108 541260 233114 541272
rect 233970 541260 233976 541272
rect 233108 541232 233976 541260
rect 233108 541220 233114 541232
rect 233970 541220 233976 541232
rect 234028 541220 234034 541272
rect 11146 540948 11152 541000
rect 11204 540988 11210 541000
rect 232038 540988 232044 541000
rect 11204 540960 232044 540988
rect 11204 540948 11210 540960
rect 232038 540948 232044 540960
rect 232096 540948 232102 541000
rect 453758 540948 453764 541000
rect 453816 540988 453822 541000
rect 462682 540988 462688 541000
rect 453816 540960 462688 540988
rect 453816 540948 453822 540960
rect 462682 540948 462688 540960
rect 462740 540948 462746 541000
rect 42794 540200 42800 540252
rect 42852 540240 42858 540252
rect 225690 540240 225696 540252
rect 42852 540212 225696 540240
rect 42852 540200 42858 540212
rect 225690 540200 225696 540212
rect 225748 540200 225754 540252
rect 223114 539588 223120 539640
rect 223172 539628 223178 539640
rect 232038 539628 232044 539640
rect 223172 539600 232044 539628
rect 223172 539588 223178 539600
rect 232038 539588 232044 539600
rect 232096 539588 232102 539640
rect 189718 538228 189724 538280
rect 189776 538268 189782 538280
rect 232038 538268 232044 538280
rect 189776 538240 232044 538268
rect 189776 538228 189782 538240
rect 232038 538228 232044 538240
rect 232096 538228 232102 538280
rect 224586 536800 224592 536852
rect 224644 536840 224650 536852
rect 232038 536840 232044 536852
rect 224644 536812 232044 536840
rect 224644 536800 224650 536812
rect 232038 536800 232044 536812
rect 232096 536800 232102 536852
rect 453758 536800 453764 536852
rect 453816 536840 453822 536852
rect 463142 536840 463148 536852
rect 453816 536812 463148 536840
rect 453816 536800 453822 536812
rect 463142 536800 463148 536812
rect 463200 536800 463206 536852
rect 479518 536800 479524 536852
rect 479576 536840 479582 536852
rect 580166 536840 580172 536852
rect 479576 536812 580172 536840
rect 479576 536800 479582 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 453942 535440 453948 535492
rect 454000 535480 454006 535492
rect 520918 535480 520924 535492
rect 454000 535452 520924 535480
rect 454000 535440 454006 535452
rect 520918 535440 520924 535452
rect 520976 535440 520982 535492
rect 80054 534080 80060 534132
rect 80112 534120 80118 534132
rect 232038 534120 232044 534132
rect 80112 534092 232044 534120
rect 80112 534080 80118 534092
rect 232038 534080 232044 534092
rect 232096 534080 232102 534132
rect 229738 532720 229744 532772
rect 229796 532760 229802 532772
rect 232314 532760 232320 532772
rect 229796 532732 232320 532760
rect 229796 532720 229802 532732
rect 232314 532720 232320 532732
rect 232372 532720 232378 532772
rect 453942 532720 453948 532772
rect 454000 532760 454006 532772
rect 461210 532760 461216 532772
rect 454000 532732 461216 532760
rect 454000 532720 454006 532732
rect 461210 532720 461216 532732
rect 461268 532720 461274 532772
rect 1394 529932 1400 529984
rect 1452 529972 1458 529984
rect 232038 529972 232044 529984
rect 1452 529944 232044 529972
rect 1452 529932 1458 529944
rect 232038 529932 232044 529944
rect 232096 529932 232102 529984
rect 96614 528572 96620 528624
rect 96672 528612 96678 528624
rect 232038 528612 232044 528624
rect 96672 528584 232044 528612
rect 96672 528572 96678 528584
rect 232038 528572 232044 528584
rect 232096 528572 232102 528624
rect 3326 527144 3332 527196
rect 3384 527184 3390 527196
rect 19978 527184 19984 527196
rect 3384 527156 19984 527184
rect 3384 527144 3390 527156
rect 19978 527144 19984 527156
rect 20036 527144 20042 527196
rect 453942 527144 453948 527196
rect 454000 527184 454006 527196
rect 471974 527184 471980 527196
rect 454000 527156 471980 527184
rect 454000 527144 454006 527156
rect 471974 527144 471980 527156
rect 472032 527144 472038 527196
rect 224678 525784 224684 525836
rect 224736 525824 224742 525836
rect 232038 525824 232044 525836
rect 224736 525796 232044 525824
rect 224736 525784 224742 525796
rect 232038 525784 232044 525796
rect 232096 525784 232102 525836
rect 453666 524696 453672 524748
rect 453724 524736 453730 524748
rect 455782 524736 455788 524748
rect 453724 524708 455788 524736
rect 453724 524696 453730 524708
rect 455782 524696 455788 524708
rect 455840 524696 455846 524748
rect 128354 524424 128360 524476
rect 128412 524464 128418 524476
rect 232038 524464 232044 524476
rect 128412 524436 232044 524464
rect 128412 524424 128418 524436
rect 232038 524424 232044 524436
rect 232096 524424 232102 524476
rect 452930 523676 452936 523728
rect 452988 523716 452994 523728
rect 453574 523716 453580 523728
rect 452988 523688 453580 523716
rect 452988 523676 452994 523688
rect 453574 523676 453580 523688
rect 453632 523676 453638 523728
rect 4154 521636 4160 521688
rect 4212 521676 4218 521688
rect 232038 521676 232044 521688
rect 4212 521648 232044 521676
rect 4212 521636 4218 521648
rect 232038 521636 232044 521648
rect 232096 521636 232102 521688
rect 453942 521636 453948 521688
rect 454000 521676 454006 521688
rect 461578 521676 461584 521688
rect 454000 521648 461584 521676
rect 454000 521636 454006 521648
rect 461578 521636 461584 521648
rect 461636 521636 461642 521688
rect 453942 520888 453948 520940
rect 454000 520928 454006 520940
rect 457162 520928 457168 520940
rect 454000 520900 457168 520928
rect 454000 520888 454006 520900
rect 457162 520888 457168 520900
rect 457220 520888 457226 520940
rect 204254 520276 204260 520328
rect 204312 520316 204318 520328
rect 232038 520316 232044 520328
rect 204312 520288 232044 520316
rect 204312 520276 204318 520288
rect 232038 520276 232044 520288
rect 232096 520276 232102 520328
rect 223206 518916 223212 518968
rect 223264 518956 223270 518968
rect 232038 518956 232044 518968
rect 223264 518928 232044 518956
rect 223264 518916 223270 518928
rect 232038 518916 232044 518928
rect 232096 518916 232102 518968
rect 453942 518916 453948 518968
rect 454000 518956 454006 518968
rect 475470 518956 475476 518968
rect 454000 518928 475476 518956
rect 454000 518916 454006 518928
rect 475470 518916 475476 518928
rect 475528 518916 475534 518968
rect 88334 516128 88340 516180
rect 88392 516168 88398 516180
rect 232038 516168 232044 516180
rect 88392 516140 232044 516168
rect 88392 516128 88398 516140
rect 232038 516128 232044 516140
rect 232096 516128 232102 516180
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 224126 514808 224132 514820
rect 3384 514780 224132 514808
rect 3384 514768 3390 514780
rect 224126 514768 224132 514780
rect 224184 514768 224190 514820
rect 453942 514768 453948 514820
rect 454000 514808 454006 514820
rect 500218 514808 500224 514820
rect 454000 514780 500224 514808
rect 454000 514768 454006 514780
rect 500218 514768 500224 514780
rect 500276 514768 500282 514820
rect 453114 514020 453120 514072
rect 453172 514060 453178 514072
rect 453574 514060 453580 514072
rect 453172 514032 453580 514060
rect 453172 514020 453178 514032
rect 453574 514020 453580 514032
rect 453632 514020 453638 514072
rect 453758 513272 453764 513324
rect 453816 513312 453822 513324
rect 465718 513312 465724 513324
rect 453816 513284 465724 513312
rect 453816 513272 453822 513284
rect 465718 513272 465724 513284
rect 465776 513272 465782 513324
rect 227162 510620 227168 510672
rect 227220 510660 227226 510672
rect 232038 510660 232044 510672
rect 227220 510632 232044 510660
rect 227220 510620 227226 510632
rect 232038 510620 232044 510632
rect 232096 510620 232102 510672
rect 541618 510620 541624 510672
rect 541676 510660 541682 510672
rect 580166 510660 580172 510672
rect 541676 510632 580172 510660
rect 541676 510620 541682 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 453758 509260 453764 509312
rect 453816 509300 453822 509312
rect 462774 509300 462780 509312
rect 453816 509272 462780 509300
rect 453816 509260 453822 509272
rect 462774 509260 462780 509272
rect 462832 509260 462838 509312
rect 228726 506472 228732 506524
rect 228784 506512 228790 506524
rect 232038 506512 232044 506524
rect 228784 506484 232044 506512
rect 228784 506472 228790 506484
rect 232038 506472 232044 506484
rect 232096 506472 232102 506524
rect 222102 505112 222108 505164
rect 222160 505152 222166 505164
rect 232038 505152 232044 505164
rect 222160 505124 232044 505152
rect 222160 505112 222166 505124
rect 232038 505112 232044 505124
rect 232096 505112 232102 505164
rect 232958 504432 232964 504484
rect 233016 504432 233022 504484
rect 232976 504280 233004 504432
rect 232958 504228 232964 504280
rect 233016 504228 233022 504280
rect 453942 503684 453948 503736
rect 454000 503724 454006 503736
rect 464246 503724 464252 503736
rect 454000 503696 464252 503724
rect 454000 503684 454006 503696
rect 464246 503684 464252 503696
rect 464304 503684 464310 503736
rect 51074 502324 51080 502376
rect 51132 502364 51138 502376
rect 232038 502364 232044 502376
rect 51132 502336 232044 502364
rect 51132 502324 51138 502336
rect 232038 502324 232044 502336
rect 232096 502324 232102 502376
rect 3234 502256 3240 502308
rect 3292 502296 3298 502308
rect 234062 502296 234068 502308
rect 3292 502268 234068 502296
rect 3292 502256 3298 502268
rect 234062 502256 234068 502268
rect 234120 502256 234126 502308
rect 220722 500964 220728 501016
rect 220780 501004 220786 501016
rect 232038 501004 232044 501016
rect 220780 500976 232044 501004
rect 220780 500964 220786 500976
rect 232038 500964 232044 500976
rect 232096 500964 232102 501016
rect 453942 499536 453948 499588
rect 454000 499576 454006 499588
rect 548518 499576 548524 499588
rect 454000 499548 548524 499576
rect 454000 499536 454006 499548
rect 548518 499536 548524 499548
rect 548576 499536 548582 499588
rect 453942 498448 453948 498500
rect 454000 498488 454006 498500
rect 457254 498488 457260 498500
rect 454000 498460 457260 498488
rect 454000 498448 454006 498460
rect 457254 498448 457260 498460
rect 457312 498448 457318 498500
rect 179414 495456 179420 495508
rect 179472 495496 179478 495508
rect 232038 495496 232044 495508
rect 179472 495468 232044 495496
rect 179472 495456 179478 495468
rect 232038 495456 232044 495468
rect 232096 495456 232102 495508
rect 453942 492600 453948 492652
rect 454000 492640 454006 492652
rect 498838 492640 498844 492652
rect 454000 492612 498844 492640
rect 454000 492600 454006 492612
rect 498838 492600 498844 492612
rect 498896 492600 498902 492652
rect 224770 488520 224776 488572
rect 224828 488560 224834 488572
rect 232038 488560 232044 488572
rect 224828 488532 232044 488560
rect 224828 488520 224834 488532
rect 232038 488520 232044 488532
rect 232096 488520 232102 488572
rect 453758 488520 453764 488572
rect 453816 488560 453822 488572
rect 464338 488560 464344 488572
rect 453816 488532 464344 488560
rect 453816 488520 453822 488532
rect 464338 488520 464344 488532
rect 464396 488520 464402 488572
rect 453942 487432 453948 487484
rect 454000 487472 454006 487484
rect 458450 487472 458456 487484
rect 454000 487444 458456 487472
rect 454000 487432 454006 487444
rect 458450 487432 458456 487444
rect 458508 487432 458514 487484
rect 230014 485800 230020 485852
rect 230072 485840 230078 485852
rect 231854 485840 231860 485852
rect 230072 485812 231860 485840
rect 230072 485800 230078 485812
rect 231854 485800 231860 485812
rect 231912 485800 231918 485852
rect 453758 485800 453764 485852
rect 453816 485840 453822 485852
rect 480898 485840 480904 485852
rect 453816 485812 480904 485840
rect 453816 485800 453822 485812
rect 480898 485800 480904 485812
rect 480956 485800 480962 485852
rect 453942 484440 453948 484492
rect 454000 484480 454006 484492
rect 458542 484480 458548 484492
rect 454000 484452 458548 484480
rect 454000 484440 454006 484452
rect 458542 484440 458548 484452
rect 458600 484440 458606 484492
rect 213822 484372 213828 484424
rect 213880 484412 213886 484424
rect 232038 484412 232044 484424
rect 213880 484384 232044 484412
rect 213880 484372 213886 484384
rect 232038 484372 232044 484384
rect 232096 484372 232102 484424
rect 471330 484372 471336 484424
rect 471388 484412 471394 484424
rect 580166 484412 580172 484424
rect 471388 484384 580172 484412
rect 471388 484372 471394 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 453206 482740 453212 482792
rect 453264 482780 453270 482792
rect 459830 482780 459836 482792
rect 453264 482752 459836 482780
rect 453264 482740 453270 482752
rect 459830 482740 459836 482752
rect 459888 482740 459894 482792
rect 222010 481652 222016 481704
rect 222068 481692 222074 481704
rect 232038 481692 232044 481704
rect 222068 481664 232044 481692
rect 222068 481652 222074 481664
rect 232038 481652 232044 481664
rect 232096 481652 232102 481704
rect 125594 480224 125600 480276
rect 125652 480264 125658 480276
rect 232038 480264 232044 480276
rect 125652 480236 232044 480264
rect 125652 480224 125658 480236
rect 232038 480224 232044 480236
rect 232096 480224 232102 480276
rect 453758 480224 453764 480276
rect 453816 480264 453822 480276
rect 542998 480264 543004 480276
rect 453816 480236 543004 480264
rect 453816 480224 453822 480236
rect 542998 480224 543004 480236
rect 543056 480224 543062 480276
rect 52454 477504 52460 477556
rect 52512 477544 52518 477556
rect 232038 477544 232044 477556
rect 52512 477516 232044 477544
rect 52512 477504 52518 477516
rect 232038 477504 232044 477516
rect 232096 477504 232102 477556
rect 453758 477504 453764 477556
rect 453816 477544 453822 477556
rect 465718 477544 465724 477556
rect 453816 477516 465724 477544
rect 453816 477504 453822 477516
rect 465718 477504 465724 477516
rect 465776 477504 465782 477556
rect 453850 476076 453856 476128
rect 453908 476116 453914 476128
rect 549898 476116 549904 476128
rect 453908 476088 549904 476116
rect 453908 476076 453914 476088
rect 549898 476076 549904 476088
rect 549956 476076 549962 476128
rect 3326 475668 3332 475720
rect 3384 475708 3390 475720
rect 8938 475708 8944 475720
rect 3384 475680 8944 475708
rect 3384 475668 3390 475680
rect 8938 475668 8944 475680
rect 8996 475668 9002 475720
rect 120074 474716 120080 474768
rect 120132 474756 120138 474768
rect 232038 474756 232044 474768
rect 120132 474728 232044 474756
rect 120132 474716 120138 474728
rect 232038 474716 232044 474728
rect 232096 474716 232102 474768
rect 453942 474716 453948 474768
rect 454000 474756 454006 474768
rect 556798 474756 556804 474768
rect 454000 474728 556804 474756
rect 454000 474716 454006 474728
rect 556798 474716 556804 474728
rect 556856 474716 556862 474768
rect 230382 473356 230388 473408
rect 230440 473396 230446 473408
rect 231854 473396 231860 473408
rect 230440 473368 231860 473396
rect 230440 473356 230446 473368
rect 231854 473356 231860 473368
rect 231912 473356 231918 473408
rect 453942 472336 453948 472388
rect 454000 472376 454006 472388
rect 458634 472376 458640 472388
rect 454000 472348 458640 472376
rect 454000 472336 454006 472348
rect 458634 472336 458640 472348
rect 458692 472336 458698 472388
rect 55214 471996 55220 472048
rect 55272 472036 55278 472048
rect 232038 472036 232044 472048
rect 55272 472008 232044 472036
rect 55272 471996 55278 472008
rect 232038 471996 232044 472008
rect 232096 471996 232102 472048
rect 453758 471248 453764 471300
rect 453816 471288 453822 471300
rect 458266 471288 458272 471300
rect 453816 471260 458272 471288
rect 453816 471248 453822 471260
rect 458266 471248 458272 471260
rect 458324 471248 458330 471300
rect 202874 470568 202880 470620
rect 202932 470608 202938 470620
rect 232038 470608 232044 470620
rect 202932 470580 232044 470608
rect 202932 470568 202938 470580
rect 232038 470568 232044 470580
rect 232096 470568 232102 470620
rect 486510 470568 486516 470620
rect 486568 470608 486574 470620
rect 579614 470608 579620 470620
rect 486568 470580 579620 470608
rect 486568 470568 486574 470580
rect 579614 470568 579620 470580
rect 579672 470568 579678 470620
rect 453942 469208 453948 469260
rect 454000 469248 454006 469260
rect 529198 469248 529204 469260
rect 454000 469220 529204 469248
rect 454000 469208 454006 469220
rect 529198 469208 529204 469220
rect 529256 469208 529262 469260
rect 452654 468528 452660 468580
rect 452712 468568 452718 468580
rect 454402 468568 454408 468580
rect 452712 468540 454408 468568
rect 452712 468528 452718 468540
rect 454402 468528 454408 468540
rect 454460 468528 454466 468580
rect 453574 466624 453580 466676
rect 453632 466664 453638 466676
rect 455966 466664 455972 466676
rect 453632 466636 455972 466664
rect 453632 466624 453638 466636
rect 455966 466624 455972 466636
rect 456024 466624 456030 466676
rect 218146 465060 218152 465112
rect 218204 465100 218210 465112
rect 232038 465100 232044 465112
rect 218204 465072 232044 465100
rect 218204 465060 218210 465072
rect 232038 465060 232044 465072
rect 232096 465060 232102 465112
rect 218238 464312 218244 464364
rect 218296 464352 218302 464364
rect 222746 464352 222752 464364
rect 218296 464324 222752 464352
rect 218296 464312 218302 464324
rect 222746 464312 222752 464324
rect 222804 464312 222810 464364
rect 453206 464176 453212 464228
rect 453264 464216 453270 464228
rect 455414 464216 455420 464228
rect 453264 464188 455420 464216
rect 453264 464176 453270 464188
rect 455414 464176 455420 464188
rect 455472 464176 455478 464228
rect 57974 463700 57980 463752
rect 58032 463740 58038 463752
rect 232038 463740 232044 463752
rect 58032 463712 232044 463740
rect 58032 463700 58038 463712
rect 232038 463700 232044 463712
rect 232096 463700 232102 463752
rect 226886 462340 226892 462392
rect 226944 462380 226950 462392
rect 232038 462380 232044 462392
rect 226944 462352 232044 462380
rect 226944 462340 226950 462352
rect 232038 462340 232044 462352
rect 232096 462340 232102 462392
rect 453942 462340 453948 462392
rect 454000 462380 454006 462392
rect 475378 462380 475384 462392
rect 454000 462352 475384 462380
rect 454000 462340 454006 462352
rect 475378 462340 475384 462352
rect 475436 462340 475442 462392
rect 48314 460912 48320 460964
rect 48372 460952 48378 460964
rect 232038 460952 232044 460964
rect 48372 460924 232044 460952
rect 48372 460912 48378 460924
rect 232038 460912 232044 460924
rect 232096 460912 232102 460964
rect 164234 459552 164240 459604
rect 164292 459592 164298 459604
rect 232038 459592 232044 459604
rect 164292 459564 232044 459592
rect 164292 459552 164298 459564
rect 232038 459552 232044 459564
rect 232096 459552 232102 459604
rect 453942 459552 453948 459604
rect 454000 459592 454006 459604
rect 504358 459592 504364 459604
rect 454000 459564 504364 459592
rect 454000 459552 454006 459564
rect 504358 459552 504364 459564
rect 504416 459552 504422 459604
rect 452654 458396 452660 458448
rect 452712 458436 452718 458448
rect 454310 458436 454316 458448
rect 452712 458408 454316 458436
rect 452712 458396 452718 458408
rect 454310 458396 454316 458408
rect 454368 458396 454374 458448
rect 220630 458192 220636 458244
rect 220688 458232 220694 458244
rect 231946 458232 231952 458244
rect 220688 458204 231952 458232
rect 220688 458192 220694 458204
rect 231946 458192 231952 458204
rect 232004 458192 232010 458244
rect 216582 456764 216588 456816
rect 216640 456804 216646 456816
rect 232038 456804 232044 456816
rect 216640 456776 232044 456804
rect 216640 456764 216646 456776
rect 232038 456764 232044 456776
rect 232096 456764 232102 456816
rect 19978 456696 19984 456748
rect 20036 456736 20042 456748
rect 231946 456736 231952 456748
rect 20036 456708 231952 456736
rect 20036 456696 20042 456708
rect 231946 456696 231952 456708
rect 232004 456696 232010 456748
rect 453666 455404 453672 455456
rect 453724 455444 453730 455456
rect 462866 455444 462872 455456
rect 453724 455416 462872 455444
rect 453724 455404 453730 455416
rect 462866 455404 462872 455416
rect 462924 455404 462930 455456
rect 453942 454248 453948 454300
rect 454000 454288 454006 454300
rect 457346 454288 457352 454300
rect 454000 454260 457352 454288
rect 454000 454248 454006 454260
rect 457346 454248 457352 454260
rect 457404 454248 457410 454300
rect 228634 454044 228640 454096
rect 228692 454084 228698 454096
rect 232038 454084 232044 454096
rect 228692 454056 232044 454084
rect 228692 454044 228698 454056
rect 232038 454044 232044 454056
rect 232096 454044 232102 454096
rect 228542 452616 228548 452668
rect 228600 452656 228606 452668
rect 232038 452656 232044 452668
rect 228600 452628 232044 452656
rect 228600 452616 228606 452628
rect 232038 452616 232044 452628
rect 232096 452616 232102 452668
rect 453942 452616 453948 452668
rect 454000 452656 454006 452668
rect 465442 452656 465448 452668
rect 454000 452628 465448 452656
rect 454000 452616 454006 452628
rect 465442 452616 465448 452628
rect 465500 452616 465506 452668
rect 153194 451256 153200 451308
rect 153252 451296 153258 451308
rect 232038 451296 232044 451308
rect 153252 451268 232044 451296
rect 153252 451256 153258 451268
rect 232038 451256 232044 451268
rect 232096 451256 232102 451308
rect 453574 450168 453580 450220
rect 453632 450208 453638 450220
rect 455874 450208 455880 450220
rect 453632 450180 455880 450208
rect 453632 450168 453638 450180
rect 455874 450168 455880 450180
rect 455932 450168 455938 450220
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 227346 449868 227352 449880
rect 3384 449840 227352 449868
rect 3384 449828 3390 449840
rect 227346 449828 227352 449840
rect 227404 449828 227410 449880
rect 453022 447448 453028 447500
rect 453080 447488 453086 447500
rect 454494 447488 454500 447500
rect 453080 447460 454500 447488
rect 453080 447448 453086 447460
rect 454494 447448 454500 447460
rect 454552 447448 454558 447500
rect 453942 444728 453948 444780
rect 454000 444768 454006 444780
rect 460014 444768 460020 444780
rect 454000 444740 460020 444768
rect 454000 444728 454006 444740
rect 460014 444728 460020 444740
rect 460072 444728 460078 444780
rect 229646 444388 229652 444440
rect 229704 444428 229710 444440
rect 232314 444428 232320 444440
rect 229704 444400 232320 444428
rect 229704 444388 229710 444400
rect 232314 444388 232320 444400
rect 232372 444388 232378 444440
rect 220538 442960 220544 443012
rect 220596 443000 220602 443012
rect 232038 443000 232044 443012
rect 220596 442972 232044 443000
rect 220596 442960 220602 442972
rect 232038 442960 232044 442972
rect 232096 442960 232102 443012
rect 225874 441600 225880 441652
rect 225932 441640 225938 441652
rect 232038 441640 232044 441652
rect 225932 441612 232044 441640
rect 225932 441600 225938 441612
rect 232038 441600 232044 441612
rect 232096 441600 232102 441652
rect 228266 440240 228272 440292
rect 228324 440280 228330 440292
rect 232038 440280 232044 440292
rect 228324 440252 232044 440280
rect 228324 440240 228330 440252
rect 232038 440240 232044 440252
rect 232096 440240 232102 440292
rect 453942 440240 453948 440292
rect 454000 440280 454006 440292
rect 544378 440280 544384 440292
rect 454000 440252 544384 440280
rect 454000 440240 454006 440252
rect 544378 440240 544384 440252
rect 544436 440240 544442 440292
rect 453850 440172 453856 440224
rect 453908 440212 453914 440224
rect 502978 440212 502984 440224
rect 453908 440184 502984 440212
rect 453908 440172 453914 440184
rect 502978 440172 502984 440184
rect 503036 440172 503042 440224
rect 453942 437452 453948 437504
rect 454000 437492 454006 437504
rect 489178 437492 489184 437504
rect 454000 437464 489184 437492
rect 454000 437452 454006 437464
rect 489178 437452 489184 437464
rect 489236 437452 489242 437504
rect 453942 436092 453948 436144
rect 454000 436132 454006 436144
rect 461302 436132 461308 436144
rect 454000 436104 461308 436132
rect 454000 436092 454006 436104
rect 461302 436092 461308 436104
rect 461360 436092 461366 436144
rect 453666 435072 453672 435124
rect 453724 435112 453730 435124
rect 456058 435112 456064 435124
rect 453724 435084 456064 435112
rect 453724 435072 453730 435084
rect 456058 435072 456064 435084
rect 456116 435072 456122 435124
rect 158714 433304 158720 433356
rect 158772 433344 158778 433356
rect 231946 433344 231952 433356
rect 158772 433316 231952 433344
rect 158772 433304 158778 433316
rect 231946 433304 231952 433316
rect 232004 433304 232010 433356
rect 79318 433236 79324 433288
rect 79376 433276 79382 433288
rect 232038 433276 232044 433288
rect 79376 433248 232044 433276
rect 79376 433236 79382 433248
rect 232038 433236 232044 433248
rect 232096 433236 232102 433288
rect 453942 430584 453948 430636
rect 454000 430624 454006 430636
rect 526438 430624 526444 430636
rect 454000 430596 526444 430624
rect 454000 430584 454006 430596
rect 526438 430584 526444 430596
rect 526496 430584 526502 430636
rect 462958 429836 462964 429888
rect 463016 429876 463022 429888
rect 580166 429876 580172 429888
rect 463016 429848 580172 429876
rect 463016 429836 463022 429848
rect 580166 429836 580172 429848
rect 580224 429836 580230 429888
rect 229554 429156 229560 429208
rect 229612 429196 229618 429208
rect 231854 429196 231860 429208
rect 229612 429168 231860 429196
rect 229612 429156 229618 429168
rect 231854 429156 231860 429168
rect 231912 429156 231918 429208
rect 91094 427796 91100 427848
rect 91152 427836 91158 427848
rect 232038 427836 232044 427848
rect 91152 427808 232044 427836
rect 91152 427796 91158 427808
rect 232038 427796 232044 427808
rect 232096 427796 232102 427848
rect 453942 427796 453948 427848
rect 454000 427836 454006 427848
rect 525058 427836 525064 427848
rect 454000 427808 525064 427836
rect 454000 427796 454006 427808
rect 525058 427796 525064 427808
rect 525116 427796 525122 427848
rect 85574 426436 85580 426488
rect 85632 426476 85638 426488
rect 232038 426476 232044 426488
rect 85632 426448 232044 426476
rect 85632 426436 85638 426448
rect 232038 426436 232044 426448
rect 232096 426436 232102 426488
rect 453942 426436 453948 426488
rect 454000 426476 454006 426488
rect 494054 426476 494060 426488
rect 454000 426448 494060 426476
rect 454000 426436 454006 426448
rect 494054 426436 494060 426448
rect 494112 426436 494118 426488
rect 168374 425076 168380 425128
rect 168432 425116 168438 425128
rect 232038 425116 232044 425128
rect 168432 425088 232044 425116
rect 168432 425076 168438 425088
rect 232038 425076 232044 425088
rect 232096 425076 232102 425128
rect 453942 425076 453948 425128
rect 454000 425116 454006 425128
rect 555418 425116 555424 425128
rect 454000 425088 555424 425116
rect 454000 425076 454006 425088
rect 555418 425076 555424 425088
rect 555476 425076 555482 425128
rect 452746 425008 452752 425060
rect 452804 425048 452810 425060
rect 541618 425048 541624 425060
rect 452804 425020 541624 425048
rect 452804 425008 452810 425020
rect 541618 425008 541624 425020
rect 541676 425008 541682 425060
rect 122834 423648 122840 423700
rect 122892 423688 122898 423700
rect 232038 423688 232044 423700
rect 122892 423660 232044 423688
rect 122892 423648 122898 423660
rect 232038 423648 232044 423660
rect 232096 423648 232102 423700
rect 3142 422288 3148 422340
rect 3200 422328 3206 422340
rect 228450 422328 228456 422340
rect 3200 422300 228456 422328
rect 3200 422288 3206 422300
rect 228450 422288 228456 422300
rect 228508 422288 228514 422340
rect 453942 420928 453948 420980
rect 454000 420968 454006 420980
rect 463878 420968 463884 420980
rect 454000 420940 463884 420968
rect 454000 420928 454006 420940
rect 463878 420928 463884 420940
rect 463936 420928 463942 420980
rect 209774 419500 209780 419552
rect 209832 419540 209838 419552
rect 232038 419540 232044 419552
rect 209832 419512 232044 419540
rect 209832 419500 209838 419512
rect 232038 419500 232044 419512
rect 232096 419500 232102 419552
rect 453666 418208 453672 418260
rect 453724 418248 453730 418260
rect 456150 418248 456156 418260
rect 453724 418220 456156 418248
rect 453724 418208 453730 418220
rect 456150 418208 456156 418220
rect 456208 418208 456214 418260
rect 491938 418140 491944 418192
rect 491996 418180 492002 418192
rect 579706 418180 579712 418192
rect 491996 418152 579712 418180
rect 491996 418140 492002 418152
rect 579706 418140 579712 418152
rect 579764 418140 579770 418192
rect 453206 416848 453212 416900
rect 453264 416888 453270 416900
rect 455506 416888 455512 416900
rect 453264 416860 455512 416888
rect 453264 416848 453270 416860
rect 455506 416848 455512 416860
rect 455564 416848 455570 416900
rect 227438 415420 227444 415472
rect 227496 415460 227502 415472
rect 231946 415460 231952 415472
rect 227496 415432 231952 415460
rect 227496 415420 227502 415432
rect 231946 415420 231952 415432
rect 232004 415420 232010 415472
rect 453942 413176 453948 413228
rect 454000 413216 454006 413228
rect 458726 413216 458732 413228
rect 454000 413188 458732 413216
rect 454000 413176 454006 413188
rect 458726 413176 458732 413188
rect 458784 413176 458790 413228
rect 227530 412632 227536 412684
rect 227588 412672 227594 412684
rect 232038 412672 232044 412684
rect 227588 412644 232044 412672
rect 227588 412632 227594 412644
rect 232038 412632 232044 412644
rect 232096 412632 232102 412684
rect 82814 409912 82820 409964
rect 82872 409952 82878 409964
rect 232038 409952 232044 409964
rect 82872 409924 232044 409952
rect 82872 409912 82878 409924
rect 232038 409912 232044 409924
rect 232096 409912 232102 409964
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 225690 409884 225696 409896
rect 3384 409856 225696 409884
rect 3384 409844 3390 409856
rect 225690 409844 225696 409856
rect 225748 409844 225754 409896
rect 452654 408824 452660 408876
rect 452712 408864 452718 408876
rect 454586 408864 454592 408876
rect 452712 408836 454592 408864
rect 452712 408824 452718 408836
rect 454586 408824 454592 408836
rect 454644 408824 454650 408876
rect 10318 408416 10324 408468
rect 10376 408456 10382 408468
rect 232038 408456 232044 408468
rect 10376 408428 232044 408456
rect 10376 408416 10382 408428
rect 232038 408416 232044 408428
rect 232096 408416 232102 408468
rect 453758 407192 453764 407244
rect 453816 407232 453822 407244
rect 456242 407232 456248 407244
rect 453816 407204 456248 407232
rect 453816 407192 453822 407204
rect 456242 407192 456248 407204
rect 456300 407192 456306 407244
rect 453942 407056 453948 407108
rect 454000 407096 454006 407108
rect 491938 407096 491944 407108
rect 454000 407068 491944 407096
rect 454000 407056 454006 407068
rect 491938 407056 491944 407068
rect 491996 407056 492002 407108
rect 453758 404880 453764 404932
rect 453816 404920 453822 404932
rect 460106 404920 460112 404932
rect 453816 404892 460112 404920
rect 453816 404880 453822 404892
rect 460106 404880 460112 404892
rect 460164 404880 460170 404932
rect 565078 404336 565084 404388
rect 565136 404376 565142 404388
rect 580166 404376 580172 404388
rect 565136 404348 580172 404376
rect 565136 404336 565142 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 132494 401616 132500 401668
rect 132552 401656 132558 401668
rect 232038 401656 232044 401668
rect 132552 401628 232044 401656
rect 132552 401616 132558 401628
rect 232038 401616 232044 401628
rect 232096 401616 232102 401668
rect 453942 401616 453948 401668
rect 454000 401656 454006 401668
rect 463050 401656 463056 401668
rect 454000 401628 463056 401656
rect 454000 401616 454006 401628
rect 463050 401616 463056 401628
rect 463108 401616 463114 401668
rect 452654 400188 452660 400240
rect 452712 400228 452718 400240
rect 454678 400228 454684 400240
rect 452712 400200 454684 400228
rect 452712 400188 452718 400200
rect 454678 400188 454684 400200
rect 454736 400188 454742 400240
rect 190454 398828 190460 398880
rect 190512 398868 190518 398880
rect 232038 398868 232044 398880
rect 190512 398840 232044 398868
rect 190512 398828 190518 398840
rect 232038 398828 232044 398840
rect 232096 398828 232102 398880
rect 453758 398828 453764 398880
rect 453816 398868 453822 398880
rect 465534 398868 465540 398880
rect 453816 398840 465540 398868
rect 453816 398828 453822 398840
rect 465534 398828 465540 398840
rect 465592 398828 465598 398880
rect 232406 398080 232412 398132
rect 232464 398120 232470 398132
rect 233142 398120 233148 398132
rect 232464 398092 233148 398120
rect 232464 398080 232470 398092
rect 233142 398080 233148 398092
rect 233200 398080 233206 398132
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 3384 397480 11008 397508
rect 3384 397468 3390 397480
rect 10980 397440 11008 397480
rect 228910 397468 228916 397520
rect 228968 397508 228974 397520
rect 232038 397508 232044 397520
rect 228968 397480 232044 397508
rect 228968 397468 228974 397480
rect 232038 397468 232044 397480
rect 232096 397468 232102 397520
rect 231946 397440 231952 397452
rect 10980 397412 231952 397440
rect 231946 397400 231952 397412
rect 232004 397400 232010 397452
rect 225782 395292 225788 395344
rect 225840 395332 225846 395344
rect 234614 395332 234620 395344
rect 225840 395304 234620 395332
rect 225840 395292 225846 395304
rect 234614 395292 234620 395304
rect 234672 395292 234678 395344
rect 95234 394680 95240 394732
rect 95292 394720 95298 394732
rect 232038 394720 232044 394732
rect 95292 394692 232044 394720
rect 95292 394680 95298 394692
rect 232038 394680 232044 394692
rect 232096 394680 232102 394732
rect 453758 394680 453764 394732
rect 453816 394720 453822 394732
rect 461486 394720 461492 394732
rect 453816 394692 461492 394720
rect 453816 394680 453822 394692
rect 461486 394680 461492 394692
rect 461544 394680 461550 394732
rect 453758 393320 453764 393372
rect 453816 393360 453822 393372
rect 464430 393360 464436 393372
rect 453816 393332 464436 393360
rect 453816 393320 453822 393332
rect 464430 393320 464436 393332
rect 464488 393320 464494 393372
rect 453942 391960 453948 392012
rect 454000 392000 454006 392012
rect 491294 392000 491300 392012
rect 454000 391972 491300 392000
rect 454000 391960 454006 391972
rect 491294 391960 491300 391972
rect 491352 391960 491358 392012
rect 191834 390532 191840 390584
rect 191892 390572 191898 390584
rect 232038 390572 232044 390584
rect 191892 390544 232044 390572
rect 191892 390532 191898 390544
rect 232038 390532 232044 390544
rect 232096 390532 232102 390584
rect 453942 389172 453948 389224
rect 454000 389212 454006 389224
rect 465626 389212 465632 389224
rect 454000 389184 465632 389212
rect 454000 389172 454006 389184
rect 465626 389172 465632 389184
rect 465684 389172 465690 389224
rect 453942 386656 453948 386708
rect 454000 386696 454006 386708
rect 457438 386696 457444 386708
rect 454000 386668 457444 386696
rect 454000 386656 454006 386668
rect 457438 386656 457444 386668
rect 457496 386656 457502 386708
rect 453942 385636 453948 385688
rect 454000 385676 454006 385688
rect 456978 385676 456984 385688
rect 454000 385648 456984 385676
rect 454000 385636 454006 385648
rect 456978 385636 456984 385648
rect 457036 385636 457042 385688
rect 24854 385024 24860 385076
rect 24912 385064 24918 385076
rect 232038 385064 232044 385076
rect 24912 385036 232044 385064
rect 24912 385024 24918 385036
rect 232038 385024 232044 385036
rect 232096 385024 232102 385076
rect 195974 383664 195980 383716
rect 196032 383704 196038 383716
rect 232038 383704 232044 383716
rect 196032 383676 232044 383704
rect 196032 383664 196038 383676
rect 232038 383664 232044 383676
rect 232096 383664 232102 383716
rect 453942 383664 453948 383716
rect 454000 383704 454006 383716
rect 502978 383704 502984 383716
rect 454000 383676 502984 383704
rect 454000 383664 454006 383676
rect 502978 383664 502984 383676
rect 503036 383664 503042 383716
rect 453206 382848 453212 382900
rect 453264 382888 453270 382900
rect 460382 382888 460388 382900
rect 453264 382860 460388 382888
rect 453264 382848 453270 382860
rect 460382 382848 460388 382860
rect 460440 382848 460446 382900
rect 230198 382236 230204 382288
rect 230256 382276 230262 382288
rect 232682 382276 232688 382288
rect 230256 382248 232688 382276
rect 230256 382236 230262 382248
rect 232682 382236 232688 382248
rect 232740 382236 232746 382288
rect 453758 378768 453764 378820
rect 453816 378808 453822 378820
rect 457530 378808 457536 378820
rect 453816 378780 457536 378808
rect 453816 378768 453822 378780
rect 457530 378768 457536 378780
rect 457588 378768 457594 378820
rect 225506 378156 225512 378208
rect 225564 378196 225570 378208
rect 232038 378196 232044 378208
rect 225564 378168 232044 378196
rect 225564 378156 225570 378168
rect 232038 378156 232044 378168
rect 232096 378156 232102 378208
rect 460290 378156 460296 378208
rect 460348 378196 460354 378208
rect 580166 378196 580172 378208
rect 460348 378168 580172 378196
rect 460348 378156 460354 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 453758 375912 453764 375964
rect 453816 375952 453822 375964
rect 458818 375952 458824 375964
rect 453816 375924 458824 375952
rect 453816 375912 453822 375924
rect 458818 375912 458824 375924
rect 458876 375912 458882 375964
rect 28994 375368 29000 375420
rect 29052 375408 29058 375420
rect 232038 375408 232044 375420
rect 29052 375380 232044 375408
rect 29052 375368 29058 375380
rect 232038 375368 232044 375380
rect 232096 375368 232102 375420
rect 230290 374144 230296 374196
rect 230348 374184 230354 374196
rect 232498 374184 232504 374196
rect 230348 374156 232504 374184
rect 230348 374144 230354 374156
rect 232498 374144 232504 374156
rect 232556 374144 232562 374196
rect 230934 374008 230940 374060
rect 230992 374048 230998 374060
rect 231854 374048 231860 374060
rect 230992 374020 231860 374048
rect 230992 374008 230998 374020
rect 231854 374008 231860 374020
rect 231912 374008 231918 374060
rect 453942 372648 453948 372700
rect 454000 372688 454006 372700
rect 456978 372688 456984 372700
rect 454000 372660 456984 372688
rect 454000 372648 454006 372660
rect 456978 372648 456984 372660
rect 457036 372648 457042 372700
rect 224494 372580 224500 372632
rect 224552 372620 224558 372632
rect 232038 372620 232044 372632
rect 224552 372592 232044 372620
rect 224552 372580 224558 372592
rect 232038 372580 232044 372592
rect 232096 372580 232102 372632
rect 223022 371220 223028 371272
rect 223080 371260 223086 371272
rect 232038 371260 232044 371272
rect 223080 371232 232044 371260
rect 223080 371220 223086 371232
rect 232038 371220 232044 371232
rect 232096 371220 232102 371272
rect 453758 371220 453764 371272
rect 453816 371260 453822 371272
rect 476758 371260 476764 371272
rect 453816 371232 476764 371260
rect 453816 371220 453822 371232
rect 476758 371220 476764 371232
rect 476816 371220 476822 371272
rect 453758 369860 453764 369912
rect 453816 369900 453822 369912
rect 534074 369900 534080 369912
rect 453816 369872 534080 369900
rect 453816 369860 453822 369872
rect 534074 369860 534080 369872
rect 534132 369860 534138 369912
rect 226242 368500 226248 368552
rect 226300 368540 226306 368552
rect 232038 368540 232044 368552
rect 226300 368512 232044 368540
rect 226300 368500 226306 368512
rect 232038 368500 232044 368512
rect 232096 368500 232102 368552
rect 453758 368500 453764 368552
rect 453816 368540 453822 368552
rect 486418 368540 486424 368552
rect 453816 368512 486424 368540
rect 453816 368500 453822 368512
rect 486418 368500 486424 368512
rect 486476 368500 486482 368552
rect 453942 367208 453948 367260
rect 454000 367248 454006 367260
rect 458910 367248 458916 367260
rect 454000 367220 458916 367248
rect 454000 367208 454006 367220
rect 458910 367208 458916 367220
rect 458968 367208 458974 367260
rect 231026 367072 231032 367124
rect 231084 367112 231090 367124
rect 231854 367112 231860 367124
rect 231084 367084 231860 367112
rect 231084 367072 231090 367084
rect 231854 367072 231860 367084
rect 231912 367072 231918 367124
rect 453942 365712 453948 365764
rect 454000 365752 454006 365764
rect 464154 365752 464160 365764
rect 454000 365724 464160 365752
rect 454000 365712 454006 365724
rect 464154 365712 464160 365724
rect 464212 365712 464218 365764
rect 453758 364420 453764 364472
rect 453816 364460 453822 364472
rect 463694 364460 463700 364472
rect 453816 364432 463700 364460
rect 453816 364420 453822 364432
rect 463694 364420 463700 364432
rect 463752 364420 463758 364472
rect 461762 364352 461768 364404
rect 461820 364392 461826 364404
rect 580166 364392 580172 364404
rect 461820 364364 580172 364392
rect 461820 364352 461826 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 194594 362924 194600 362976
rect 194652 362964 194658 362976
rect 232038 362964 232044 362976
rect 194652 362936 232044 362964
rect 194652 362924 194658 362936
rect 232038 362924 232044 362936
rect 232096 362924 232102 362976
rect 227346 361564 227352 361616
rect 227404 361604 227410 361616
rect 232038 361604 232044 361616
rect 227404 361576 232044 361604
rect 227404 361564 227410 361576
rect 232038 361564 232044 361576
rect 232096 361564 232102 361616
rect 453942 361564 453948 361616
rect 454000 361604 454006 361616
rect 462314 361604 462320 361616
rect 454000 361576 462320 361604
rect 454000 361564 454006 361576
rect 462314 361564 462320 361576
rect 462372 361564 462378 361616
rect 232222 360544 232228 360596
rect 232280 360584 232286 360596
rect 233878 360584 233884 360596
rect 232280 360556 233884 360584
rect 232280 360544 232286 360556
rect 233878 360544 233884 360556
rect 233936 360544 233942 360596
rect 453942 358776 453948 358828
rect 454000 358816 454006 358828
rect 562318 358816 562324 358828
rect 454000 358788 562324 358816
rect 454000 358776 454006 358788
rect 562318 358776 562324 358788
rect 562376 358776 562382 358828
rect 453942 357484 453948 357536
rect 454000 357524 454006 357536
rect 456794 357524 456800 357536
rect 454000 357496 456800 357524
rect 454000 357484 454006 357496
rect 456794 357484 456800 357496
rect 456852 357484 456858 357536
rect 213914 356056 213920 356108
rect 213972 356096 213978 356108
rect 232038 356096 232044 356108
rect 213972 356068 232044 356096
rect 213972 356056 213978 356068
rect 232038 356056 232044 356068
rect 232096 356056 232102 356108
rect 453482 355988 453488 356040
rect 453540 356028 453546 356040
rect 459738 356028 459744 356040
rect 453540 356000 459744 356028
rect 453540 355988 453546 356000
rect 459738 355988 459744 356000
rect 459796 355988 459802 356040
rect 224402 355308 224408 355360
rect 224460 355348 224466 355360
rect 232590 355348 232596 355360
rect 224460 355320 232596 355348
rect 224460 355308 224466 355320
rect 232590 355308 232596 355320
rect 232648 355308 232654 355360
rect 451918 355104 451924 355156
rect 451976 355144 451982 355156
rect 452930 355144 452936 355156
rect 451976 355116 452936 355144
rect 451976 355104 451982 355116
rect 452930 355104 452936 355116
rect 452988 355104 452994 355156
rect 228818 351908 228824 351960
rect 228876 351948 228882 351960
rect 232038 351948 232044 351960
rect 228876 351920 232044 351948
rect 228876 351908 228882 351920
rect 232038 351908 232044 351920
rect 232096 351908 232102 351960
rect 229002 350548 229008 350600
rect 229060 350588 229066 350600
rect 232038 350588 232044 350600
rect 229060 350560 232044 350588
rect 229060 350548 229066 350560
rect 232038 350548 232044 350560
rect 232096 350548 232102 350600
rect 453390 350344 453396 350396
rect 453448 350384 453454 350396
rect 454954 350384 454960 350396
rect 453448 350356 454960 350384
rect 453448 350344 453454 350356
rect 454954 350344 454960 350356
rect 455012 350344 455018 350396
rect 232498 349800 232504 349852
rect 232556 349840 232562 349852
rect 232958 349840 232964 349852
rect 232556 349812 232964 349840
rect 232556 349800 232562 349812
rect 232958 349800 232964 349812
rect 233016 349800 233022 349852
rect 227254 349392 227260 349444
rect 227312 349432 227318 349444
rect 228358 349432 228364 349444
rect 227312 349404 228364 349432
rect 227312 349392 227318 349404
rect 228358 349392 228364 349404
rect 228416 349392 228422 349444
rect 69014 349120 69020 349172
rect 69072 349160 69078 349172
rect 232038 349160 232044 349172
rect 69072 349132 232044 349160
rect 69072 349120 69078 349132
rect 232038 349120 232044 349132
rect 232096 349120 232102 349172
rect 452562 348780 452568 348832
rect 452620 348820 452626 348832
rect 454034 348820 454040 348832
rect 452620 348792 454040 348820
rect 452620 348780 452626 348792
rect 454034 348780 454040 348792
rect 454092 348780 454098 348832
rect 228358 347760 228364 347812
rect 228416 347800 228422 347812
rect 232038 347800 232044 347812
rect 228416 347772 232044 347800
rect 228416 347760 228422 347772
rect 232038 347760 232044 347772
rect 232096 347760 232102 347812
rect 453942 347760 453948 347812
rect 454000 347800 454006 347812
rect 478874 347800 478880 347812
rect 454000 347772 478880 347800
rect 454000 347760 454006 347772
rect 478874 347760 478880 347772
rect 478932 347760 478938 347812
rect 453298 347692 453304 347744
rect 453356 347732 453362 347744
rect 454034 347732 454040 347744
rect 453356 347704 454040 347732
rect 453356 347692 453362 347704
rect 454034 347692 454040 347704
rect 454092 347692 454098 347744
rect 453942 347556 453948 347608
rect 454000 347596 454006 347608
rect 459646 347596 459652 347608
rect 454000 347568 459652 347596
rect 454000 347556 454006 347568
rect 459646 347556 459652 347568
rect 459704 347556 459710 347608
rect 230106 346400 230112 346452
rect 230164 346440 230170 346452
rect 232590 346440 232596 346452
rect 230164 346412 232596 346440
rect 230164 346400 230170 346412
rect 232590 346400 232596 346412
rect 232648 346400 232654 346452
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 59998 346372 60004 346384
rect 3384 346344 60004 346372
rect 3384 346332 3390 346344
rect 59998 346332 60004 346344
rect 60056 346332 60062 346384
rect 222930 345040 222936 345092
rect 222988 345080 222994 345092
rect 232038 345080 232044 345092
rect 222988 345052 232044 345080
rect 222988 345040 222994 345052
rect 232038 345040 232044 345052
rect 232096 345040 232102 345092
rect 201494 344972 201500 345024
rect 201552 345012 201558 345024
rect 231946 345012 231952 345024
rect 201552 344984 231952 345012
rect 201552 344972 201558 344984
rect 231946 344972 231952 344984
rect 232004 344972 232010 345024
rect 71774 344292 71780 344344
rect 71832 344332 71838 344344
rect 222746 344332 222752 344344
rect 71832 344304 222752 344332
rect 71832 344292 71838 344304
rect 222746 344292 222752 344304
rect 222804 344292 222810 344344
rect 452930 343884 452936 343936
rect 452988 343924 452994 343936
rect 454862 343924 454868 343936
rect 452988 343896 454868 343924
rect 452988 343884 452994 343896
rect 454862 343884 454868 343896
rect 454920 343884 454926 343936
rect 452378 342320 452384 342372
rect 452436 342360 452442 342372
rect 454954 342360 454960 342372
rect 452436 342332 454960 342360
rect 452436 342320 452442 342332
rect 454954 342320 454960 342332
rect 455012 342320 455018 342372
rect 102134 342252 102140 342304
rect 102192 342292 102198 342304
rect 232038 342292 232044 342304
rect 102192 342264 232044 342292
rect 102192 342252 102198 342264
rect 232038 342252 232044 342264
rect 232096 342252 232102 342304
rect 453942 342252 453948 342304
rect 454000 342292 454006 342304
rect 471238 342292 471244 342304
rect 454000 342264 471244 342292
rect 454000 342252 454006 342264
rect 471238 342252 471244 342264
rect 471296 342252 471302 342304
rect 453942 342048 453948 342100
rect 454000 342088 454006 342100
rect 458174 342088 458180 342100
rect 454000 342060 458180 342088
rect 454000 342048 454006 342060
rect 458174 342048 458180 342060
rect 458232 342048 458238 342100
rect 74534 340892 74540 340944
rect 74592 340932 74598 340944
rect 231946 340932 231952 340944
rect 74592 340904 231952 340932
rect 74592 340892 74598 340904
rect 231946 340892 231952 340904
rect 232004 340892 232010 340944
rect 21358 340824 21364 340876
rect 21416 340864 21422 340876
rect 232038 340864 232044 340876
rect 21416 340836 232044 340864
rect 21416 340824 21422 340836
rect 232038 340824 232044 340836
rect 232096 340824 232102 340876
rect 234062 338172 234068 338224
rect 234120 338212 234126 338224
rect 235994 338212 236000 338224
rect 234120 338184 236000 338212
rect 234120 338172 234126 338184
rect 235994 338172 236000 338184
rect 236052 338172 236058 338224
rect 447134 338172 447140 338224
rect 447192 338212 447198 338224
rect 465626 338212 465632 338224
rect 447192 338184 465632 338212
rect 447192 338172 447198 338184
rect 465626 338172 465632 338184
rect 465684 338172 465690 338224
rect 34514 338104 34520 338156
rect 34572 338144 34578 338156
rect 232038 338144 232044 338156
rect 34572 338116 232044 338144
rect 34572 338104 34578 338116
rect 232038 338104 232044 338116
rect 232096 338104 232102 338156
rect 226242 338036 226248 338088
rect 226300 338076 226306 338088
rect 580442 338076 580448 338088
rect 226300 338048 580448 338076
rect 226300 338036 226306 338048
rect 580442 338036 580448 338048
rect 580500 338036 580506 338088
rect 229002 337968 229008 338020
rect 229060 338008 229066 338020
rect 580534 338008 580540 338020
rect 229060 337980 580540 338008
rect 229060 337968 229066 337980
rect 580534 337968 580540 337980
rect 580592 337968 580598 338020
rect 409874 337900 409880 337952
rect 409932 337940 409938 337952
rect 452194 337940 452200 337952
rect 409932 337912 452200 337940
rect 409932 337900 409938 337912
rect 452194 337900 452200 337912
rect 452252 337900 452258 337952
rect 419534 337832 419540 337884
rect 419592 337872 419598 337884
rect 464062 337872 464068 337884
rect 419592 337844 464068 337872
rect 419592 337832 419598 337844
rect 464062 337832 464068 337844
rect 464120 337832 464126 337884
rect 405734 337764 405740 337816
rect 405792 337804 405798 337816
rect 462774 337804 462780 337816
rect 405792 337776 462780 337804
rect 405792 337764 405798 337776
rect 462774 337764 462780 337776
rect 462832 337764 462838 337816
rect 394694 337696 394700 337748
rect 394752 337736 394758 337748
rect 456794 337736 456800 337748
rect 394752 337708 456800 337736
rect 394752 337696 394758 337708
rect 456794 337696 456800 337708
rect 456852 337696 456858 337748
rect 231578 337628 231584 337680
rect 231636 337668 231642 337680
rect 244274 337668 244280 337680
rect 231636 337640 244280 337668
rect 231636 337628 231642 337640
rect 244274 337628 244280 337640
rect 244332 337628 244338 337680
rect 387794 337628 387800 337680
rect 387852 337668 387858 337680
rect 458726 337668 458732 337680
rect 387852 337640 458732 337668
rect 387852 337628 387858 337640
rect 458726 337628 458732 337640
rect 458784 337628 458790 337680
rect 225966 337560 225972 337612
rect 226024 337600 226030 337612
rect 253934 337600 253940 337612
rect 226024 337572 253940 337600
rect 226024 337560 226030 337572
rect 253934 337560 253940 337572
rect 253992 337560 253998 337612
rect 376754 337560 376760 337612
rect 376812 337600 376818 337612
rect 454126 337600 454132 337612
rect 376812 337572 454132 337600
rect 376812 337560 376818 337572
rect 454126 337560 454132 337572
rect 454184 337560 454190 337612
rect 233142 337492 233148 337544
rect 233200 337532 233206 337544
rect 262214 337532 262220 337544
rect 233200 337504 262220 337532
rect 233200 337492 233206 337504
rect 262214 337492 262220 337504
rect 262272 337492 262278 337544
rect 333974 337492 333980 337544
rect 334032 337532 334038 337544
rect 452010 337532 452016 337544
rect 334032 337504 452016 337532
rect 334032 337492 334038 337504
rect 452010 337492 452016 337504
rect 452068 337492 452074 337544
rect 233602 337424 233608 337476
rect 233660 337464 233666 337476
rect 278774 337464 278780 337476
rect 233660 337436 278780 337464
rect 233660 337424 233666 337436
rect 278774 337424 278780 337436
rect 278832 337424 278838 337476
rect 448514 337424 448520 337476
rect 448572 337464 448578 337476
rect 580626 337464 580632 337476
rect 448572 337436 580632 337464
rect 448572 337424 448578 337436
rect 580626 337424 580632 337436
rect 580684 337424 580690 337476
rect 224310 337356 224316 337408
rect 224368 337396 224374 337408
rect 243078 337396 243084 337408
rect 224368 337368 243084 337396
rect 224368 337356 224374 337368
rect 243078 337356 243084 337368
rect 243136 337356 243142 337408
rect 249794 337356 249800 337408
rect 249852 337396 249858 337408
rect 454678 337396 454684 337408
rect 249852 337368 454684 337396
rect 249852 337356 249858 337368
rect 454678 337356 454684 337368
rect 454736 337356 454742 337408
rect 427998 337288 428004 337340
rect 428056 337328 428062 337340
rect 465350 337328 465356 337340
rect 428056 337300 465356 337328
rect 428056 337288 428062 337300
rect 465350 337288 465356 337300
rect 465408 337288 465414 337340
rect 430574 337220 430580 337272
rect 430632 337260 430638 337272
rect 462866 337260 462872 337272
rect 430632 337232 462872 337260
rect 430632 337220 430638 337232
rect 462866 337220 462872 337232
rect 462924 337220 462930 337272
rect 434714 337152 434720 337204
rect 434772 337192 434778 337204
rect 455690 337192 455696 337204
rect 434772 337164 455696 337192
rect 434772 337152 434778 337164
rect 455690 337152 455696 337164
rect 455748 337152 455754 337204
rect 451274 337084 451280 337136
rect 451332 337124 451338 337136
rect 464246 337124 464252 337136
rect 451332 337096 464252 337124
rect 451332 337084 451338 337096
rect 464246 337084 464252 337096
rect 464304 337084 464310 337136
rect 227070 336812 227076 336864
rect 227128 336852 227134 336864
rect 245010 336852 245016 336864
rect 227128 336824 245016 336852
rect 227128 336812 227134 336824
rect 245010 336812 245016 336824
rect 245068 336812 245074 336864
rect 3510 336744 3516 336796
rect 3568 336784 3574 336796
rect 262398 336784 262404 336796
rect 3568 336756 262404 336784
rect 3568 336744 3574 336756
rect 262398 336744 262404 336756
rect 262456 336744 262462 336796
rect 449084 336756 450584 336784
rect 225782 336676 225788 336728
rect 225840 336716 225846 336728
rect 378318 336716 378324 336728
rect 225840 336688 378324 336716
rect 225840 336676 225846 336688
rect 378318 336676 378324 336688
rect 378376 336676 378382 336728
rect 378778 336676 378784 336728
rect 378836 336716 378842 336728
rect 380894 336716 380900 336728
rect 378836 336688 380900 336716
rect 378836 336676 378842 336688
rect 380894 336676 380900 336688
rect 380952 336676 380958 336728
rect 400858 336676 400864 336728
rect 400916 336716 400922 336728
rect 402146 336716 402152 336728
rect 400916 336688 402152 336716
rect 400916 336676 400922 336688
rect 402146 336676 402152 336688
rect 402204 336676 402210 336728
rect 422938 336676 422944 336728
rect 422996 336716 423002 336728
rect 423674 336716 423680 336728
rect 422996 336688 423680 336716
rect 422996 336676 423002 336688
rect 423674 336676 423680 336688
rect 423732 336676 423738 336728
rect 427078 336676 427084 336728
rect 427136 336716 427142 336728
rect 427906 336716 427912 336728
rect 427136 336688 427912 336716
rect 427136 336676 427142 336688
rect 427906 336676 427912 336688
rect 427964 336676 427970 336728
rect 446582 336676 446588 336728
rect 446640 336716 446646 336728
rect 449084 336716 449112 336756
rect 446640 336688 449112 336716
rect 446640 336676 446646 336688
rect 449158 336676 449164 336728
rect 449216 336716 449222 336728
rect 450446 336716 450452 336728
rect 449216 336688 450452 336716
rect 449216 336676 449222 336688
rect 450446 336676 450452 336688
rect 450504 336676 450510 336728
rect 450556 336716 450584 336756
rect 485038 336716 485044 336728
rect 450556 336688 485044 336716
rect 485038 336676 485044 336688
rect 485096 336676 485102 336728
rect 222562 336608 222568 336660
rect 222620 336648 222626 336660
rect 266354 336648 266360 336660
rect 222620 336620 266360 336648
rect 222620 336608 222626 336620
rect 266354 336608 266360 336620
rect 266412 336608 266418 336660
rect 342898 336608 342904 336660
rect 342956 336648 342962 336660
rect 461762 336648 461768 336660
rect 342956 336620 461768 336648
rect 342956 336608 342962 336620
rect 461762 336608 461768 336620
rect 461820 336608 461826 336660
rect 222746 336540 222752 336592
rect 222804 336580 222810 336592
rect 241146 336580 241152 336592
rect 222804 336552 241152 336580
rect 222804 336540 222810 336552
rect 241146 336540 241152 336552
rect 241204 336540 241210 336592
rect 244918 336540 244924 336592
rect 244976 336580 244982 336592
rect 246298 336580 246304 336592
rect 244976 336552 246304 336580
rect 244976 336540 244982 336552
rect 246298 336540 246304 336552
rect 246356 336540 246362 336592
rect 275370 336540 275376 336592
rect 275428 336580 275434 336592
rect 283650 336580 283656 336592
rect 275428 336552 283656 336580
rect 275428 336540 275434 336552
rect 283650 336540 283656 336552
rect 283708 336540 283714 336592
rect 367094 336540 367100 336592
rect 367152 336580 367158 336592
rect 464430 336580 464436 336592
rect 367152 336552 464436 336580
rect 367152 336540 367158 336552
rect 464430 336540 464436 336552
rect 464488 336540 464494 336592
rect 232406 336472 232412 336524
rect 232464 336512 232470 336524
rect 291194 336512 291200 336524
rect 232464 336484 291200 336512
rect 232464 336472 232470 336484
rect 291194 336472 291200 336484
rect 291252 336472 291258 336524
rect 357434 336472 357440 336524
rect 357492 336512 357498 336524
rect 461394 336512 461400 336524
rect 357492 336484 461400 336512
rect 357492 336472 357498 336484
rect 461394 336472 461400 336484
rect 461452 336472 461458 336524
rect 229830 336404 229836 336456
rect 229888 336444 229894 336456
rect 296714 336444 296720 336456
rect 229888 336416 296720 336444
rect 229888 336404 229894 336416
rect 296714 336404 296720 336416
rect 296772 336404 296778 336456
rect 441338 336404 441344 336456
rect 441396 336444 441402 336456
rect 462958 336444 462964 336456
rect 441396 336416 462964 336444
rect 441396 336404 441402 336416
rect 462958 336404 462964 336416
rect 463016 336404 463022 336456
rect 224954 336336 224960 336388
rect 225012 336376 225018 336388
rect 460014 336376 460020 336388
rect 225012 336348 460020 336376
rect 225012 336336 225018 336348
rect 460014 336336 460020 336348
rect 460072 336336 460078 336388
rect 21358 336268 21364 336320
rect 21416 336308 21422 336320
rect 269114 336308 269120 336320
rect 21416 336280 269120 336308
rect 21416 336268 21422 336280
rect 269114 336268 269120 336280
rect 269172 336268 269178 336320
rect 277394 336268 277400 336320
rect 277452 336308 277458 336320
rect 454586 336308 454592 336320
rect 277452 336280 454592 336308
rect 277452 336268 277458 336280
rect 454586 336268 454592 336280
rect 454644 336268 454650 336320
rect 165614 336200 165620 336252
rect 165672 336240 165678 336252
rect 463050 336240 463056 336252
rect 165672 336212 463056 336240
rect 165672 336200 165678 336212
rect 463050 336200 463056 336212
rect 463108 336200 463114 336252
rect 24118 336132 24124 336184
rect 24176 336172 24182 336184
rect 323578 336172 323584 336184
rect 24176 336144 323584 336172
rect 24176 336132 24182 336144
rect 323578 336132 323584 336144
rect 323636 336132 323642 336184
rect 342254 336132 342260 336184
rect 342312 336172 342318 336184
rect 459922 336172 459928 336184
rect 342312 336144 459928 336172
rect 342312 336132 342318 336144
rect 459922 336132 459928 336144
rect 459980 336132 459986 336184
rect 28258 336064 28264 336116
rect 28316 336104 28322 336116
rect 413094 336104 413100 336116
rect 28316 336076 413100 336104
rect 28316 336064 28322 336076
rect 413094 336064 413100 336076
rect 413152 336064 413158 336116
rect 424962 336064 424968 336116
rect 425020 336104 425026 336116
rect 486510 336104 486516 336116
rect 425020 336076 486516 336104
rect 425020 336064 425026 336076
rect 486510 336064 486516 336076
rect 486568 336064 486574 336116
rect 26878 335996 26884 336048
rect 26936 336036 26942 336048
rect 416958 336036 416964 336048
rect 26936 336008 416964 336036
rect 26936 335996 26942 336008
rect 416958 335996 416964 336008
rect 417016 335996 417022 336048
rect 420178 335996 420184 336048
rect 420236 336036 420242 336048
rect 436738 336036 436744 336048
rect 420236 336008 436744 336036
rect 420236 335996 420242 336008
rect 436738 335996 436744 336008
rect 436796 335996 436802 336048
rect 440234 335996 440240 336048
rect 440292 336036 440298 336048
rect 457254 336036 457260 336048
rect 440292 336008 457260 336036
rect 440292 335996 440298 336008
rect 457254 335996 457260 336008
rect 457312 335996 457318 336048
rect 222838 335928 222844 335980
rect 222896 335968 222902 335980
rect 233234 335968 233240 335980
rect 222896 335940 233240 335968
rect 222896 335928 222902 335940
rect 233234 335928 233240 335940
rect 233292 335928 233298 335980
rect 280798 335928 280804 335980
rect 280856 335968 280862 335980
rect 282362 335968 282368 335980
rect 280856 335940 282368 335968
rect 280856 335928 280862 335940
rect 282362 335928 282368 335940
rect 282420 335928 282426 335980
rect 381538 335928 381544 335980
rect 381596 335968 381602 335980
rect 389266 335968 389272 335980
rect 381596 335940 389272 335968
rect 381596 335928 381602 335940
rect 389266 335928 389272 335940
rect 389324 335928 389330 335980
rect 405366 335928 405372 335980
rect 405424 335968 405430 335980
rect 448514 335968 448520 335980
rect 405424 335940 448520 335968
rect 405424 335928 405430 335940
rect 448514 335928 448520 335940
rect 448572 335928 448578 335980
rect 225690 335860 225696 335912
rect 225748 335900 225754 335912
rect 234890 335900 234896 335912
rect 225748 335872 234896 335900
rect 225748 335860 225754 335872
rect 234890 335860 234896 335872
rect 234948 335860 234954 335912
rect 407114 335860 407120 335912
rect 407172 335900 407178 335912
rect 433334 335900 433340 335912
rect 407172 335872 433340 335900
rect 407172 335860 407178 335872
rect 433334 335860 433340 335872
rect 433392 335860 433398 335912
rect 404998 335792 405004 335844
rect 405056 335832 405062 335844
rect 425974 335832 425980 335844
rect 405056 335804 425980 335832
rect 405056 335792 405062 335804
rect 425974 335792 425980 335804
rect 426032 335792 426038 335844
rect 320174 335656 320180 335708
rect 320232 335696 320238 335708
rect 451826 335696 451832 335708
rect 320232 335668 451832 335696
rect 320232 335656 320238 335668
rect 451826 335656 451832 335668
rect 451884 335656 451890 335708
rect 360930 335588 360936 335640
rect 360988 335628 360994 335640
rect 366082 335628 366088 335640
rect 360988 335600 366088 335628
rect 360988 335588 360994 335600
rect 366082 335588 366088 335600
rect 366140 335588 366146 335640
rect 380986 335588 380992 335640
rect 381044 335628 381050 335640
rect 456886 335628 456892 335640
rect 381044 335600 456892 335628
rect 381044 335588 381050 335600
rect 456886 335588 456892 335600
rect 456944 335588 456950 335640
rect 232866 334908 232872 334960
rect 232924 334948 232930 334960
rect 282914 334948 282920 334960
rect 232924 334920 282920 334948
rect 232924 334908 232930 334920
rect 282914 334908 282920 334920
rect 282972 334908 282978 334960
rect 364334 334908 364340 334960
rect 364392 334948 364398 334960
rect 455966 334948 455972 334960
rect 364392 334920 455972 334948
rect 364392 334908 364398 334920
rect 455966 334908 455972 334920
rect 456024 334908 456030 334960
rect 233970 334840 233976 334892
rect 234028 334880 234034 334892
rect 298094 334880 298100 334892
rect 234028 334852 298100 334880
rect 234028 334840 234034 334852
rect 298094 334840 298100 334852
rect 298152 334840 298158 334892
rect 340874 334840 340880 334892
rect 340932 334880 340938 334892
rect 452102 334880 452108 334892
rect 340932 334852 452108 334880
rect 340932 334840 340938 334852
rect 452102 334840 452108 334852
rect 452160 334840 452166 334892
rect 230934 334772 230940 334824
rect 230992 334812 230998 334824
rect 375374 334812 375380 334824
rect 230992 334784 375380 334812
rect 230992 334772 230998 334784
rect 375374 334772 375380 334784
rect 375432 334772 375438 334824
rect 415394 334772 415400 334824
rect 415452 334812 415458 334824
rect 451734 334812 451740 334824
rect 415452 334784 451740 334812
rect 415452 334772 415458 334784
rect 451734 334772 451740 334784
rect 451792 334772 451798 334824
rect 234614 334704 234620 334756
rect 234672 334744 234678 334756
rect 241514 334744 241520 334756
rect 234672 334716 241520 334744
rect 234672 334704 234678 334716
rect 241514 334704 241520 334716
rect 241572 334704 241578 334756
rect 259638 334704 259644 334756
rect 259696 334744 259702 334756
rect 452654 334744 452660 334756
rect 259696 334716 452660 334744
rect 259696 334704 259702 334716
rect 452654 334704 452660 334716
rect 452712 334704 452718 334756
rect 232130 334636 232136 334688
rect 232188 334676 232194 334688
rect 438854 334676 438860 334688
rect 232188 334648 438860 334676
rect 232188 334636 232194 334648
rect 438854 334636 438860 334648
rect 438912 334636 438918 334688
rect 44174 334568 44180 334620
rect 44232 334608 44238 334620
rect 453482 334608 453488 334620
rect 44232 334580 453488 334608
rect 44232 334568 44238 334580
rect 453482 334568 453488 334580
rect 453540 334568 453546 334620
rect 23474 333888 23480 333940
rect 23532 333928 23538 333940
rect 324866 333928 324872 333940
rect 23532 333900 324872 333928
rect 23532 333888 23538 333900
rect 324866 333888 324872 333900
rect 324924 333888 324930 333940
rect 398742 333888 398748 333940
rect 398800 333928 398806 333940
rect 565078 333928 565084 333940
rect 398800 333900 565084 333928
rect 398800 333888 398806 333900
rect 565078 333888 565084 333900
rect 565136 333888 565142 333940
rect 286870 333820 286876 333872
rect 286928 333860 286934 333872
rect 471330 333860 471336 333872
rect 286928 333832 471336 333860
rect 286928 333820 286934 333832
rect 471330 333820 471336 333832
rect 471388 333820 471394 333872
rect 131758 333752 131764 333804
rect 131816 333792 131822 333804
rect 397270 333792 397276 333804
rect 131816 333764 397276 333792
rect 131816 333752 131822 333764
rect 397270 333752 397276 333764
rect 397328 333752 397334 333804
rect 418154 333752 418160 333804
rect 418212 333792 418218 333804
rect 462682 333792 462688 333804
rect 418212 333764 462688 333792
rect 418212 333752 418218 333764
rect 462682 333752 462688 333764
rect 462740 333752 462746 333804
rect 255222 333684 255228 333736
rect 255280 333724 255286 333736
rect 477494 333724 477500 333736
rect 255280 333696 477500 333724
rect 255280 333684 255286 333696
rect 477494 333684 477500 333696
rect 477552 333684 477558 333736
rect 253382 333616 253388 333668
rect 253440 333656 253446 333668
rect 460290 333656 460296 333668
rect 253440 333628 460296 333656
rect 253440 333616 253446 333628
rect 460290 333616 460296 333628
rect 460348 333616 460354 333668
rect 275278 333548 275284 333600
rect 275336 333588 275342 333600
rect 479518 333588 479524 333600
rect 275336 333560 479524 333588
rect 275336 333548 275342 333560
rect 479518 333548 479524 333560
rect 479576 333548 479582 333600
rect 157978 333480 157984 333532
rect 158036 333520 158042 333532
rect 356054 333520 356060 333532
rect 158036 333492 356060 333520
rect 158036 333480 158042 333492
rect 356054 333480 356060 333492
rect 356112 333480 356118 333532
rect 373994 333480 374000 333532
rect 374052 333520 374058 333532
rect 451642 333520 451648 333532
rect 374052 333492 451648 333520
rect 374052 333480 374058 333492
rect 451642 333480 451648 333492
rect 451700 333480 451706 333532
rect 225506 333412 225512 333464
rect 225564 333452 225570 333464
rect 231854 333452 231860 333464
rect 225564 333424 231860 333452
rect 225564 333412 225570 333424
rect 231854 333412 231860 333424
rect 231912 333412 231918 333464
rect 248414 333412 248420 333464
rect 248472 333452 248478 333464
rect 465258 333452 465264 333464
rect 248472 333424 465264 333452
rect 248472 333412 248478 333424
rect 465258 333412 465264 333424
rect 465316 333412 465322 333464
rect 201494 333344 201500 333396
rect 201552 333384 201558 333396
rect 457438 333384 457444 333396
rect 201552 333356 457444 333384
rect 201552 333344 201558 333356
rect 457438 333344 457444 333356
rect 457496 333344 457502 333396
rect 200114 333276 200120 333328
rect 200172 333316 200178 333328
rect 462314 333316 462320 333328
rect 200172 333288 462320 333316
rect 200172 333276 200178 333288
rect 462314 333276 462320 333288
rect 462372 333276 462378 333328
rect 129734 333208 129740 333260
rect 129792 333248 129798 333260
rect 458174 333248 458180 333260
rect 129792 333220 458180 333248
rect 129792 333208 129798 333220
rect 458174 333208 458180 333220
rect 458232 333208 458238 333260
rect 224126 333140 224132 333192
rect 224184 333180 224190 333192
rect 390554 333180 390560 333192
rect 224184 333152 390560 333180
rect 224184 333140 224190 333152
rect 390554 333140 390560 333152
rect 390612 333140 390618 333192
rect 429194 333140 429200 333192
rect 429252 333180 429258 333192
rect 463694 333180 463700 333192
rect 429252 333152 463700 333180
rect 429252 333140 429258 333152
rect 463694 333140 463700 333152
rect 463752 333140 463758 333192
rect 40034 333072 40040 333124
rect 40092 333112 40098 333124
rect 311986 333112 311992 333124
rect 40092 333084 311992 333112
rect 40092 333072 40098 333084
rect 311986 333072 311992 333084
rect 312044 333072 312050 333124
rect 347774 333072 347780 333124
rect 347832 333112 347838 333124
rect 452286 333112 452292 333124
rect 347832 333084 452292 333112
rect 347832 333072 347838 333084
rect 452286 333072 452292 333084
rect 452344 333072 452350 333124
rect 352006 333004 352012 333056
rect 352064 333044 352070 333056
rect 451550 333044 451556 333056
rect 352064 333016 451556 333044
rect 352064 333004 352070 333016
rect 451550 333004 451556 333016
rect 451608 333004 451614 333056
rect 234798 331984 234804 332036
rect 234856 332024 234862 332036
rect 271874 332024 271880 332036
rect 234856 331996 271880 332024
rect 234856 331984 234862 331996
rect 271874 331984 271880 331996
rect 271932 331984 271938 332036
rect 232774 331916 232780 331968
rect 232832 331956 232838 331968
rect 303614 331956 303620 331968
rect 232832 331928 303620 331956
rect 232832 331916 232838 331928
rect 303614 331916 303620 331928
rect 303672 331916 303678 331968
rect 307754 331916 307760 331968
rect 307812 331956 307818 331968
rect 456242 331956 456248 331968
rect 307812 331928 456248 331956
rect 307812 331916 307818 331928
rect 456242 331916 456248 331928
rect 456300 331916 456306 331968
rect 267826 331848 267832 331900
rect 267884 331888 267890 331900
rect 453022 331888 453028 331900
rect 267884 331860 453028 331888
rect 267884 331848 267890 331860
rect 453022 331848 453028 331860
rect 453080 331848 453086 331900
rect 231302 330624 231308 330676
rect 231360 330664 231366 330676
rect 317506 330664 317512 330676
rect 231360 330636 317512 330664
rect 231360 330624 231366 330636
rect 317506 330624 317512 330636
rect 317564 330624 317570 330676
rect 349154 330624 349160 330676
rect 349212 330664 349218 330676
rect 454494 330664 454500 330676
rect 349212 330636 454500 330664
rect 349212 330624 349218 330636
rect 454494 330624 454500 330636
rect 454552 330624 454558 330676
rect 233694 330556 233700 330608
rect 233752 330596 233758 330608
rect 281534 330596 281540 330608
rect 233752 330568 281540 330596
rect 233752 330556 233758 330568
rect 281534 330556 281540 330568
rect 281592 330556 281598 330608
rect 311894 330556 311900 330608
rect 311952 330596 311958 330608
rect 455782 330596 455788 330608
rect 311952 330568 455788 330596
rect 311952 330556 311958 330568
rect 455782 330556 455788 330568
rect 455840 330556 455846 330608
rect 231670 330488 231676 330540
rect 231728 330528 231734 330540
rect 382274 330528 382280 330540
rect 231728 330500 382280 330528
rect 231728 330488 231734 330500
rect 382274 330488 382280 330500
rect 382332 330488 382338 330540
rect 270586 330420 270592 330472
rect 270644 330460 270650 330472
rect 271414 330460 271420 330472
rect 270644 330432 271420 330460
rect 270644 330420 270650 330432
rect 271414 330420 271420 330432
rect 271472 330420 271478 330472
rect 346394 330420 346400 330472
rect 346452 330460 346458 330472
rect 347406 330460 347412 330472
rect 346452 330432 347412 330460
rect 346452 330420 346458 330432
rect 347406 330420 347412 330432
rect 347464 330420 347470 330472
rect 228910 329060 228916 329112
rect 228968 329100 228974 329112
rect 400214 329100 400220 329112
rect 228968 329072 400220 329100
rect 228968 329060 228974 329072
rect 400214 329060 400220 329072
rect 400272 329060 400278 329112
rect 284294 327768 284300 327820
rect 284352 327808 284358 327820
rect 455598 327808 455604 327820
rect 284352 327780 455604 327808
rect 284352 327768 284358 327780
rect 455598 327768 455604 327780
rect 455656 327768 455662 327820
rect 183554 327700 183560 327752
rect 183612 327740 183618 327752
rect 454402 327740 454408 327752
rect 183612 327712 454408 327740
rect 183612 327700 183618 327712
rect 454402 327700 454408 327712
rect 454460 327700 454466 327752
rect 394786 326748 394792 326800
rect 394844 326788 394850 326800
rect 395706 326788 395712 326800
rect 394844 326760 395712 326788
rect 394844 326748 394850 326760
rect 395706 326748 395712 326760
rect 395764 326748 395770 326800
rect 233878 326476 233884 326528
rect 233936 326516 233942 326528
rect 383654 326516 383660 326528
rect 233936 326488 383660 326516
rect 233936 326476 233942 326488
rect 383654 326476 383660 326488
rect 383712 326476 383718 326528
rect 251174 326408 251180 326460
rect 251232 326448 251238 326460
rect 453758 326448 453764 326460
rect 251232 326420 453764 326448
rect 251232 326408 251238 326420
rect 453758 326408 453764 326420
rect 453816 326408 453822 326460
rect 223574 326340 223580 326392
rect 223632 326380 223638 326392
rect 456150 326380 456156 326392
rect 223632 326352 456156 326380
rect 223632 326340 223638 326352
rect 456150 326340 456156 326352
rect 456208 326340 456214 326392
rect 329834 325592 329840 325644
rect 329892 325632 329898 325644
rect 580166 325632 580172 325644
rect 329892 325604 580172 325632
rect 329892 325592 329898 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 231394 325116 231400 325168
rect 231452 325156 231458 325168
rect 353294 325156 353300 325168
rect 231452 325128 353300 325156
rect 231452 325116 231458 325128
rect 353294 325116 353300 325128
rect 353352 325116 353358 325168
rect 229646 325048 229652 325100
rect 229704 325088 229710 325100
rect 477494 325088 477500 325100
rect 229704 325060 477500 325088
rect 229704 325048 229710 325060
rect 477494 325048 477500 325060
rect 477552 325048 477558 325100
rect 184934 324980 184940 325032
rect 184992 325020 184998 325032
rect 449894 325020 449900 325032
rect 184992 324992 449900 325020
rect 184992 324980 184998 324992
rect 449894 324980 449900 324992
rect 449952 324980 449958 325032
rect 121454 324912 121460 324964
rect 121512 324952 121518 324964
rect 457346 324952 457352 324964
rect 121512 324924 457352 324952
rect 121512 324912 121518 324924
rect 457346 324912 457352 324924
rect 457404 324912 457410 324964
rect 233786 323620 233792 323672
rect 233844 323660 233850 323672
rect 346486 323660 346492 323672
rect 233844 323632 346492 323660
rect 233844 323620 233850 323632
rect 346486 323620 346492 323632
rect 346544 323620 346550 323672
rect 228542 323552 228548 323604
rect 228600 323592 228606 323604
rect 280154 323592 280160 323604
rect 228600 323564 280160 323592
rect 228600 323552 228606 323564
rect 280154 323552 280160 323564
rect 280212 323552 280218 323604
rect 292574 323552 292580 323604
rect 292632 323592 292638 323604
rect 454218 323592 454224 323604
rect 292632 323564 454224 323592
rect 292632 323552 292638 323564
rect 454218 323552 454224 323564
rect 454276 323552 454282 323604
rect 340966 322260 340972 322312
rect 341024 322300 341030 322312
rect 457162 322300 457168 322312
rect 341024 322272 457168 322300
rect 341024 322260 341030 322272
rect 457162 322260 457168 322272
rect 457220 322260 457226 322312
rect 81434 322192 81440 322244
rect 81492 322232 81498 322244
rect 225690 322232 225696 322244
rect 81492 322204 225696 322232
rect 81492 322192 81498 322204
rect 225690 322192 225696 322204
rect 225748 322192 225754 322244
rect 229738 322192 229744 322244
rect 229796 322232 229802 322244
rect 420914 322232 420920 322244
rect 229796 322204 420920 322232
rect 229796 322192 229802 322204
rect 420914 322192 420920 322204
rect 420972 322192 420978 322244
rect 231118 320832 231124 320884
rect 231176 320872 231182 320884
rect 510614 320872 510620 320884
rect 231176 320844 510620 320872
rect 231176 320832 231182 320844
rect 510614 320832 510620 320844
rect 510672 320832 510678 320884
rect 3510 320084 3516 320136
rect 3568 320124 3574 320136
rect 220170 320124 220176 320136
rect 3568 320096 220176 320124
rect 3568 320084 3574 320096
rect 220170 320084 220176 320096
rect 220228 320084 220234 320136
rect 231026 319540 231032 319592
rect 231084 319580 231090 319592
rect 310514 319580 310520 319592
rect 231084 319552 310520 319580
rect 231084 319540 231090 319552
rect 310514 319540 310520 319552
rect 310572 319540 310578 319592
rect 229554 319472 229560 319524
rect 229612 319512 229618 319524
rect 393406 319512 393412 319524
rect 229612 319484 393412 319512
rect 229612 319472 229618 319484
rect 393406 319472 393412 319484
rect 393464 319472 393470 319524
rect 78674 319404 78680 319456
rect 78732 319444 78738 319456
rect 453206 319444 453212 319456
rect 78732 319416 453212 319444
rect 78732 319404 78738 319416
rect 453206 319404 453212 319416
rect 453264 319404 453270 319456
rect 228634 318044 228640 318096
rect 228692 318084 228698 318096
rect 276014 318084 276020 318096
rect 228692 318056 276020 318084
rect 228692 318044 228698 318056
rect 276014 318044 276020 318056
rect 276072 318044 276078 318096
rect 284386 318044 284392 318096
rect 284444 318084 284450 318096
rect 454310 318084 454316 318096
rect 284444 318056 454316 318084
rect 284444 318044 284450 318056
rect 454310 318044 454316 318056
rect 454368 318044 454374 318096
rect 387242 316684 387248 316736
rect 387300 316724 387306 316736
rect 568574 316724 568580 316736
rect 387300 316696 568580 316724
rect 387300 316684 387306 316696
rect 568574 316684 568580 316696
rect 568632 316684 568638 316736
rect 260834 315324 260840 315376
rect 260892 315364 260898 315376
rect 449158 315364 449164 315376
rect 260892 315336 449164 315364
rect 260892 315324 260898 315336
rect 449158 315324 449164 315336
rect 449216 315324 449222 315376
rect 189074 315256 189080 315308
rect 189132 315296 189138 315308
rect 448514 315296 448520 315308
rect 189132 315268 448520 315296
rect 189132 315256 189138 315268
rect 448514 315256 448520 315268
rect 448572 315256 448578 315308
rect 556798 313216 556804 313268
rect 556856 313256 556862 313268
rect 580166 313256 580172 313268
rect 556856 313228 580172 313256
rect 556856 313216 556862 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 49694 312536 49700 312588
rect 49752 312576 49758 312588
rect 458634 312576 458640 312588
rect 49752 312548 458640 312576
rect 49752 312536 49758 312548
rect 458634 312536 458640 312548
rect 458692 312536 458698 312588
rect 345014 309816 345020 309868
rect 345072 309856 345078 309868
rect 437474 309856 437480 309868
rect 345072 309828 437480 309856
rect 345072 309816 345078 309828
rect 437474 309816 437480 309828
rect 437532 309816 437538 309868
rect 329834 309748 329840 309800
rect 329892 309788 329898 309800
rect 457622 309788 457628 309800
rect 329892 309760 457628 309788
rect 329892 309748 329898 309760
rect 457622 309748 457628 309760
rect 457680 309748 457686 309800
rect 369854 308456 369860 308508
rect 369912 308496 369918 308508
rect 436094 308496 436100 308508
rect 369912 308468 436100 308496
rect 369912 308456 369918 308468
rect 436094 308456 436100 308468
rect 436152 308456 436158 308508
rect 198734 308388 198740 308440
rect 198792 308428 198798 308440
rect 453114 308428 453120 308440
rect 198792 308400 453120 308428
rect 198792 308388 198798 308400
rect 453114 308388 453120 308400
rect 453172 308388 453178 308440
rect 216674 307028 216680 307080
rect 216732 307068 216738 307080
rect 456058 307068 456064 307080
rect 216732 307040 456064 307068
rect 216732 307028 216738 307040
rect 456058 307028 456064 307040
rect 456116 307028 456122 307080
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 317598 306320 317604 306332
rect 3568 306292 317604 306320
rect 3568 306280 3574 306292
rect 317598 306280 317604 306292
rect 317656 306280 317662 306332
rect 324314 305668 324320 305720
rect 324372 305708 324378 305720
rect 374086 305708 374092 305720
rect 324372 305680 374092 305708
rect 324372 305668 324378 305680
rect 374086 305668 374092 305680
rect 374144 305668 374150 305720
rect 389174 305668 389180 305720
rect 389232 305708 389238 305720
rect 400306 305708 400312 305720
rect 389232 305680 400312 305708
rect 389232 305668 389238 305680
rect 400306 305668 400312 305680
rect 400364 305668 400370 305720
rect 433426 305668 433432 305720
rect 433484 305708 433490 305720
rect 547874 305708 547880 305720
rect 433484 305680 547880 305708
rect 433484 305668 433490 305680
rect 547874 305668 547880 305680
rect 547932 305668 547938 305720
rect 234154 305600 234160 305652
rect 234212 305640 234218 305652
rect 498194 305640 498200 305652
rect 234212 305612 498200 305640
rect 234212 305600 234218 305612
rect 498194 305600 498200 305612
rect 498252 305600 498258 305652
rect 345106 303016 345112 303068
rect 345164 303056 345170 303068
rect 402974 303056 402980 303068
rect 345164 303028 402980 303056
rect 345164 303016 345170 303028
rect 402974 303016 402980 303028
rect 403032 303016 403038 303068
rect 150434 302948 150440 303000
rect 150492 302988 150498 303000
rect 346578 302988 346584 303000
rect 150492 302960 346584 302988
rect 150492 302948 150498 302960
rect 346578 302948 346584 302960
rect 346636 302948 346642 303000
rect 394878 302948 394884 303000
rect 394936 302988 394942 303000
rect 533338 302988 533344 303000
rect 394936 302960 533344 302988
rect 394936 302948 394942 302960
rect 533338 302948 533344 302960
rect 533396 302948 533402 303000
rect 115934 302880 115940 302932
rect 115992 302920 115998 302932
rect 458542 302920 458548 302932
rect 115992 302892 458548 302920
rect 115992 302880 115998 302892
rect 458542 302880 458548 302892
rect 458600 302880 458606 302932
rect 234338 301452 234344 301504
rect 234396 301492 234402 301504
rect 580626 301492 580632 301504
rect 234396 301464 580632 301492
rect 234396 301452 234402 301464
rect 580626 301452 580632 301464
rect 580684 301452 580690 301504
rect 103514 300160 103520 300212
rect 103572 300200 103578 300212
rect 259546 300200 259552 300212
rect 103572 300172 259552 300200
rect 103572 300160 103578 300172
rect 259546 300160 259552 300172
rect 259604 300160 259610 300212
rect 232682 300092 232688 300144
rect 232740 300132 232746 300144
rect 408586 300132 408592 300144
rect 232740 300104 408592 300132
rect 232740 300092 232746 300104
rect 408586 300092 408592 300104
rect 408644 300092 408650 300144
rect 468570 299412 468576 299464
rect 468628 299452 468634 299464
rect 580166 299452 580172 299464
rect 468628 299424 580172 299452
rect 468628 299412 468634 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 173894 297372 173900 297424
rect 173952 297412 173958 297424
rect 455874 297412 455880 297424
rect 173952 297384 455880 297412
rect 173952 297372 173958 297384
rect 455874 297372 455880 297384
rect 455932 297372 455938 297424
rect 228726 296012 228732 296064
rect 228784 296052 228790 296064
rect 322934 296052 322940 296064
rect 228784 296024 322940 296052
rect 228784 296012 228790 296024
rect 322934 296012 322940 296024
rect 322992 296012 322998 296064
rect 309134 295944 309140 295996
rect 309192 295984 309198 295996
rect 484394 295984 484400 295996
rect 309192 295956 484400 295984
rect 309192 295944 309198 295956
rect 484394 295944 484400 295956
rect 484452 295944 484458 295996
rect 284478 294652 284484 294704
rect 284536 294692 284542 294704
rect 502334 294692 502340 294704
rect 284536 294664 502340 294692
rect 284536 294652 284542 294664
rect 502334 294652 502340 294664
rect 502392 294652 502398 294704
rect 84194 294584 84200 294636
rect 84252 294624 84258 294636
rect 458450 294624 458456 294636
rect 84252 294596 458456 294624
rect 84252 294584 84258 294596
rect 458450 294584 458456 294596
rect 458508 294584 458514 294636
rect 3510 293904 3516 293956
rect 3568 293944 3574 293956
rect 461210 293944 461216 293956
rect 3568 293916 461216 293944
rect 3568 293904 3574 293916
rect 461210 293904 461216 293916
rect 461268 293904 461274 293956
rect 231486 291864 231492 291916
rect 231544 291904 231550 291916
rect 335446 291904 335452 291916
rect 231544 291876 335452 291904
rect 231544 291864 231550 291876
rect 335446 291864 335452 291876
rect 335504 291864 335510 291916
rect 9674 291796 9680 291848
rect 9732 291836 9738 291848
rect 251266 291836 251272 291848
rect 9732 291808 251272 291836
rect 9732 291796 9738 291808
rect 251266 291796 251272 291808
rect 251324 291796 251330 291848
rect 320266 291796 320272 291848
rect 320324 291836 320330 291848
rect 556246 291836 556252 291848
rect 320324 291808 556252 291836
rect 320324 291796 320330 291808
rect 556246 291796 556252 291808
rect 556304 291796 556310 291848
rect 59354 290504 59360 290556
rect 59412 290544 59418 290556
rect 242986 290544 242992 290556
rect 59412 290516 242992 290544
rect 59412 290504 59418 290516
rect 242986 290504 242992 290516
rect 243044 290504 243050 290556
rect 231210 290436 231216 290488
rect 231268 290476 231274 290488
rect 516134 290476 516140 290488
rect 231268 290448 516140 290476
rect 231268 290436 231274 290448
rect 516134 290436 516140 290448
rect 516192 290436 516198 290488
rect 172514 289076 172520 289128
rect 172572 289116 172578 289128
rect 438946 289116 438952 289128
rect 172572 289088 438952 289116
rect 172572 289076 172578 289088
rect 438946 289076 438952 289088
rect 439004 289076 439010 289128
rect 147674 284928 147680 284980
rect 147732 284968 147738 284980
rect 341058 284968 341064 284980
rect 147732 284940 341064 284968
rect 147732 284928 147738 284940
rect 341058 284928 341064 284940
rect 341116 284928 341122 284980
rect 361574 284928 361580 284980
rect 361632 284968 361638 284980
rect 549254 284968 549260 284980
rect 361632 284940 549260 284968
rect 361632 284928 361638 284940
rect 549254 284928 549260 284940
rect 549312 284928 549318 284980
rect 316126 282140 316132 282192
rect 316184 282180 316190 282192
rect 378134 282180 378140 282192
rect 316184 282152 378140 282180
rect 316184 282140 316190 282152
rect 378134 282140 378140 282152
rect 378192 282140 378198 282192
rect 144914 280780 144920 280832
rect 144972 280820 144978 280832
rect 280246 280820 280252 280832
rect 144972 280792 280252 280820
rect 144972 280780 144978 280792
rect 280246 280780 280252 280792
rect 280304 280780 280310 280832
rect 292666 280780 292672 280832
rect 292724 280820 292730 280832
rect 396074 280820 396080 280832
rect 292724 280792 396080 280820
rect 292724 280780 292730 280792
rect 396074 280780 396080 280792
rect 396132 280780 396138 280832
rect 234522 273164 234528 273216
rect 234580 273204 234586 273216
rect 580166 273204 580172 273216
rect 234580 273176 580172 273204
rect 234580 273164 234586 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 53834 272484 53840 272536
rect 53892 272524 53898 272536
rect 255314 272524 255320 272536
rect 53892 272496 255320 272524
rect 53892 272484 53898 272496
rect 255314 272484 255320 272496
rect 255372 272484 255378 272536
rect 313274 272484 313280 272536
rect 313332 272524 313338 272536
rect 567838 272524 567844 272536
rect 313332 272496 567844 272524
rect 313332 272484 313338 272496
rect 567838 272484 567844 272496
rect 567896 272484 567902 272536
rect 226334 269764 226340 269816
rect 226392 269804 226398 269816
rect 385126 269804 385132 269816
rect 226392 269776 385132 269804
rect 226392 269764 226398 269776
rect 385126 269764 385132 269776
rect 385184 269764 385190 269816
rect 369946 268404 369952 268456
rect 370004 268444 370010 268456
rect 467834 268444 467840 268456
rect 370004 268416 467840 268444
rect 370004 268404 370010 268416
rect 467834 268404 467840 268416
rect 467892 268404 467898 268456
rect 135346 268336 135352 268388
rect 135404 268376 135410 268388
rect 375466 268376 375472 268388
rect 135404 268348 375472 268376
rect 135404 268336 135410 268348
rect 375466 268336 375472 268348
rect 375524 268336 375530 268388
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 461486 267696 461492 267708
rect 3568 267668 461492 267696
rect 3568 267656 3574 267668
rect 461486 267656 461492 267668
rect 461544 267656 461550 267708
rect 294046 262964 294052 263016
rect 294104 263004 294110 263016
rect 427078 263004 427084 263016
rect 294104 262976 427084 263004
rect 294104 262964 294110 262976
rect 427078 262964 427084 262976
rect 427136 262964 427142 263016
rect 142154 262828 142160 262880
rect 142212 262868 142218 262880
rect 293954 262868 293960 262880
rect 142212 262840 293960 262868
rect 142212 262828 142218 262840
rect 293954 262828 293960 262840
rect 294012 262828 294018 262880
rect 151814 257320 151820 257372
rect 151872 257360 151878 257372
rect 328454 257360 328460 257372
rect 151872 257332 328460 257360
rect 151872 257320 151878 257332
rect 328454 257320 328460 257332
rect 328512 257320 328518 257372
rect 227162 255960 227168 256012
rect 227220 256000 227226 256012
rect 411254 256000 411260 256012
rect 227220 255972 411260 256000
rect 227220 255960 227226 255972
rect 411254 255960 411260 255972
rect 411312 255960 411318 256012
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 459830 255252 459836 255264
rect 3200 255224 459836 255252
rect 3200 255212 3206 255224
rect 459830 255212 459836 255224
rect 459888 255212 459894 255264
rect 226886 254532 226892 254584
rect 226944 254572 226950 254584
rect 422386 254572 422392 254584
rect 226944 254544 422392 254572
rect 226944 254532 226950 254544
rect 422386 254532 422392 254544
rect 422444 254532 422450 254584
rect 89714 250452 89720 250504
rect 89772 250492 89778 250504
rect 422938 250492 422944 250504
rect 89772 250464 422944 250492
rect 89772 250452 89778 250464
rect 422938 250452 422944 250464
rect 422996 250452 423002 250504
rect 100754 247664 100760 247716
rect 100812 247704 100818 247716
rect 360194 247704 360200 247716
rect 100812 247676 360200 247704
rect 100812 247664 100818 247676
rect 360194 247664 360200 247676
rect 360252 247664 360258 247716
rect 33134 246304 33140 246356
rect 33192 246344 33198 246356
rect 306374 246344 306380 246356
rect 33192 246316 306380 246344
rect 33192 246304 33198 246316
rect 306374 246304 306380 246316
rect 306432 246304 306438 246356
rect 225874 245556 225880 245608
rect 225932 245596 225938 245608
rect 580166 245596 580172 245608
rect 225932 245568 580172 245596
rect 225932 245556 225938 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 66254 239368 66260 239420
rect 66312 239408 66318 239420
rect 458266 239408 458272 239420
rect 66312 239380 458272 239408
rect 66312 239368 66318 239380
rect 458266 239368 458272 239380
rect 458324 239368 458330 239420
rect 70394 235220 70400 235272
rect 70452 235260 70458 235272
rect 382458 235260 382464 235272
rect 70452 235232 382464 235260
rect 70452 235220 70458 235232
rect 382458 235220 382464 235232
rect 382516 235220 382522 235272
rect 230014 233928 230020 233980
rect 230072 233968 230078 233980
rect 386414 233968 386420 233980
rect 230072 233940 386420 233968
rect 230072 233928 230078 233940
rect 386414 233928 386420 233940
rect 386472 233928 386478 233980
rect 13814 233860 13820 233912
rect 13872 233900 13878 233912
rect 405826 233900 405832 233912
rect 13872 233872 405832 233900
rect 13872 233860 13878 233872
rect 405826 233860 405832 233872
rect 405884 233860 405890 233912
rect 99374 232500 99380 232552
rect 99432 232540 99438 232552
rect 278866 232540 278872 232552
rect 99432 232512 278872 232540
rect 99432 232500 99438 232512
rect 278866 232500 278872 232512
rect 278924 232500 278930 232552
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 447226 215268 447232 215280
rect 3384 215240 447232 215268
rect 3384 215228 3390 215240
rect 447226 215228 447232 215240
rect 447284 215228 447290 215280
rect 376846 206932 376852 206984
rect 376904 206972 376910 206984
rect 579982 206972 579988 206984
rect 376904 206944 579988 206972
rect 376904 206932 376910 206944
rect 579982 206932 579988 206944
rect 580040 206932 580046 206984
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 461302 202824 461308 202836
rect 3476 202796 461308 202824
rect 3476 202784 3482 202796
rect 461302 202784 461308 202796
rect 461360 202784 461366 202836
rect 475470 193128 475476 193180
rect 475528 193168 475534 193180
rect 580166 193168 580172 193180
rect 475528 193140 580172 193168
rect 475528 193128 475534 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 464154 189020 464160 189032
rect 3476 188992 464160 189020
rect 3476 188980 3482 188992
rect 464154 188980 464160 188992
rect 464212 188980 464218 189032
rect 208394 180072 208400 180124
rect 208452 180112 208458 180124
rect 452838 180112 452844 180124
rect 208452 180084 452844 180112
rect 208452 180072 208458 180084
rect 452838 180072 452844 180084
rect 452896 180072 452902 180124
rect 247034 179324 247040 179376
rect 247092 179364 247098 179376
rect 580166 179364 580172 179376
rect 247092 179336 580172 179364
rect 247092 179324 247098 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 169754 174496 169760 174548
rect 169812 174536 169818 174548
rect 455506 174536 455512 174548
rect 169812 174508 455512 174536
rect 169812 174496 169818 174508
rect 455506 174496 455512 174508
rect 455564 174496 455570 174548
rect 233050 173136 233056 173188
rect 233108 173176 233114 173188
rect 423674 173176 423680 173188
rect 233108 173148 423680 173176
rect 233108 173136 233114 173148
rect 423674 173136 423680 173148
rect 423732 173136 423738 173188
rect 224586 166948 224592 167000
rect 224644 166988 224650 167000
rect 580166 166988 580172 167000
rect 224644 166960 580172 166988
rect 224644 166948 224650 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 211154 164840 211160 164892
rect 211212 164880 211218 164892
rect 431954 164880 431960 164892
rect 211212 164852 431960 164880
rect 211212 164840 211218 164852
rect 431954 164840 431960 164852
rect 432012 164840 432018 164892
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 211798 164200 211804 164212
rect 3292 164172 211804 164200
rect 3292 164160 3298 164172
rect 211798 164160 211804 164172
rect 211856 164160 211862 164212
rect 35986 157972 35992 158024
rect 36044 158012 36050 158024
rect 244918 158012 244924 158024
rect 36044 157984 244924 158012
rect 36044 157972 36050 157984
rect 244918 157972 244924 157984
rect 244976 157972 244982 158024
rect 527818 153144 527824 153196
rect 527876 153184 527882 153196
rect 579982 153184 579988 153196
rect 527876 153156 579988 153184
rect 527876 153144 527882 153156
rect 579982 153144 579988 153156
rect 580040 153144 580046 153196
rect 300854 152464 300860 152516
rect 300912 152504 300918 152516
rect 527174 152504 527180 152516
rect 300912 152476 527180 152504
rect 300912 152464 300918 152476
rect 527174 152464 527180 152476
rect 527232 152464 527238 152516
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 385034 150396 385040 150408
rect 3476 150368 385040 150396
rect 3476 150356 3482 150368
rect 385034 150356 385040 150368
rect 385092 150356 385098 150408
rect 62114 145528 62120 145580
rect 62172 145568 62178 145580
rect 275278 145568 275284 145580
rect 62172 145540 275284 145568
rect 62172 145528 62178 145540
rect 275278 145528 275284 145540
rect 275336 145528 275342 145580
rect 287054 139340 287060 139392
rect 287112 139380 287118 139392
rect 580166 139380 580172 139392
rect 287112 139352 580172 139380
rect 287112 139340 287118 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 469858 138660 469864 138712
rect 469916 138700 469922 138712
rect 580258 138700 580264 138712
rect 469916 138672 580264 138700
rect 469916 138660 469922 138672
rect 580258 138660 580264 138672
rect 580316 138660 580322 138712
rect 263594 123428 263600 123480
rect 263652 123468 263658 123480
rect 331306 123468 331312 123480
rect 263652 123440 331312 123468
rect 263652 123428 263658 123440
rect 331306 123428 331312 123440
rect 331364 123428 331370 123480
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 206278 111772 206284 111784
rect 3476 111744 206284 111772
rect 3476 111732 3482 111744
rect 206278 111732 206284 111744
rect 206336 111732 206342 111784
rect 480898 100648 480904 100700
rect 480956 100688 480962 100700
rect 580166 100688 580172 100700
rect 480956 100660 580172 100688
rect 480956 100648 480962 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 267918 97968 267924 97980
rect 3476 97940 267924 97968
rect 3476 97928 3482 97940
rect 267918 97928 267924 97940
rect 267976 97928 267982 97980
rect 295334 91740 295340 91792
rect 295392 91780 295398 91792
rect 474734 91780 474740 91792
rect 295392 91752 474740 91780
rect 295392 91740 295398 91752
rect 474734 91740 474740 91752
rect 474792 91740 474798 91792
rect 30374 90312 30380 90364
rect 30432 90352 30438 90364
rect 343634 90352 343640 90364
rect 30432 90324 343640 90352
rect 30432 90312 30438 90324
rect 343634 90312 343640 90324
rect 343692 90312 343698 90364
rect 209866 87592 209872 87644
rect 209924 87632 209930 87644
rect 452746 87632 452752 87644
rect 209924 87604 452752 87632
rect 209924 87592 209930 87604
rect 452746 87592 452752 87604
rect 452804 87592 452810 87644
rect 224678 86912 224684 86964
rect 224736 86952 224742 86964
rect 580166 86952 580172 86964
rect 224736 86924 580172 86952
rect 224736 86912 224742 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 231762 86232 231768 86284
rect 231820 86272 231826 86284
rect 365714 86272 365720 86284
rect 231820 86244 365720 86272
rect 231820 86232 231826 86244
rect 365714 86232 365720 86244
rect 365772 86232 365778 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 199378 85524 199384 85536
rect 3200 85496 199384 85524
rect 3200 85484 3206 85496
rect 199378 85484 199384 85496
rect 199436 85484 199442 85536
rect 232314 80656 232320 80708
rect 232372 80696 232378 80708
rect 416774 80696 416780 80708
rect 232372 80668 416780 80696
rect 232372 80656 232378 80668
rect 416774 80656 416780 80668
rect 416832 80656 416838 80708
rect 223114 73108 223120 73160
rect 223172 73148 223178 73160
rect 580166 73148 580172 73160
rect 223172 73120 580172 73148
rect 223172 73108 223178 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 200758 71720 200764 71732
rect 3476 71692 200764 71720
rect 3476 71680 3482 71692
rect 200758 71680 200764 71692
rect 200816 71680 200822 71732
rect 77294 69640 77300 69692
rect 77352 69680 77358 69692
rect 378778 69680 378784 69692
rect 77352 69652 378784 69680
rect 77352 69640 77358 69652
rect 378778 69640 378784 69652
rect 378836 69640 378842 69692
rect 85666 65492 85672 65544
rect 85724 65532 85730 65544
rect 360838 65532 360844 65544
rect 85724 65504 360844 65532
rect 85724 65492 85730 65504
rect 360838 65492 360844 65504
rect 360896 65492 360902 65544
rect 69106 64132 69112 64184
rect 69164 64172 69170 64184
rect 383746 64172 383752 64184
rect 69164 64144 383752 64172
rect 69164 64132 69170 64144
rect 383746 64132 383752 64144
rect 383804 64132 383810 64184
rect 227438 59984 227444 60036
rect 227496 60024 227502 60036
rect 397454 60024 397460 60036
rect 227496 59996 397460 60024
rect 227496 59984 227502 59996
rect 397454 59984 397460 59996
rect 397512 59984 397518 60036
rect 241606 57196 241612 57248
rect 241664 57236 241670 57248
rect 368566 57236 368572 57248
rect 241664 57208 368572 57236
rect 241664 57196 241670 57208
rect 368566 57196 368572 57208
rect 368624 57196 368630 57248
rect 149054 55836 149060 55888
rect 149112 55876 149118 55888
rect 404998 55876 405004 55888
rect 149112 55848 405004 55876
rect 149112 55836 149118 55848
rect 404998 55836 405004 55848
rect 405056 55836 405062 55888
rect 287054 54476 287060 54528
rect 287112 54516 287118 54528
rect 434806 54516 434812 54528
rect 287112 54488 434812 54516
rect 287112 54476 287118 54488
rect 434806 54476 434812 54488
rect 434864 54476 434870 54528
rect 27614 51756 27620 51808
rect 27672 51796 27678 51808
rect 269298 51796 269304 51808
rect 27672 51768 269304 51796
rect 27672 51756 27678 51768
rect 269298 51756 269304 51768
rect 269356 51756 269362 51808
rect 269206 51688 269212 51740
rect 269264 51728 269270 51740
rect 400858 51728 400864 51740
rect 269264 51700 400864 51728
rect 269264 51688 269270 51700
rect 400858 51688 400864 51700
rect 400916 51688 400922 51740
rect 321554 47608 321560 47660
rect 321612 47648 321618 47660
rect 528554 47648 528560 47660
rect 321612 47620 528560 47648
rect 321612 47608 321618 47620
rect 528554 47608 528560 47620
rect 528612 47608 528618 47660
rect 234614 47540 234620 47592
rect 234672 47580 234678 47592
rect 455414 47580 455420 47592
rect 234672 47552 455420 47580
rect 234672 47540 234678 47552
rect 455414 47540 455420 47552
rect 455472 47540 455478 47592
rect 507118 46860 507124 46912
rect 507176 46900 507182 46912
rect 580166 46900 580172 46912
rect 507176 46872 580172 46900
rect 507176 46860 507182 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 334066 46180 334072 46232
rect 334124 46220 334130 46232
rect 489914 46220 489920 46232
rect 334124 46192 489920 46220
rect 334124 46180 334130 46192
rect 489914 46180 489920 46192
rect 489972 46180 489978 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 338114 45540 338120 45552
rect 3476 45512 338120 45540
rect 3476 45500 3482 45512
rect 338114 45500 338120 45512
rect 338172 45500 338178 45552
rect 298186 43392 298192 43444
rect 298244 43432 298250 43444
rect 470594 43432 470600 43444
rect 298244 43404 470600 43432
rect 298244 43392 298250 43404
rect 470594 43392 470600 43404
rect 470652 43392 470658 43444
rect 398926 39312 398932 39364
rect 398984 39352 398990 39364
rect 459646 39352 459652 39364
rect 398984 39324 459652 39352
rect 398984 39312 398990 39324
rect 459646 39312 459652 39324
rect 459704 39312 459710 39364
rect 40034 35164 40040 35216
rect 40092 35204 40098 35216
rect 453666 35204 453672 35216
rect 40092 35176 453672 35204
rect 40092 35164 40098 35176
rect 453666 35164 453672 35176
rect 453724 35164 453730 35216
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 456978 33096 456984 33108
rect 3568 33068 456984 33096
rect 3568 33056 3574 33068
rect 456978 33056 456984 33068
rect 457036 33056 457042 33108
rect 473998 33056 474004 33108
rect 474056 33096 474062 33108
rect 580166 33096 580172 33108
rect 474056 33068 580172 33096
rect 474056 33056 474062 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 237466 32376 237472 32428
rect 237524 32416 237530 32428
rect 372706 32416 372712 32428
rect 237524 32388 372712 32416
rect 237524 32376 237530 32388
rect 372706 32376 372712 32388
rect 372764 32376 372770 32428
rect 228266 31016 228272 31068
rect 228324 31056 228330 31068
rect 332686 31056 332692 31068
rect 228324 31028 332692 31056
rect 228324 31016 228330 31028
rect 332686 31016 332692 31028
rect 332744 31016 332750 31068
rect 489178 31016 489184 31068
rect 489236 31056 489242 31068
rect 506474 31056 506480 31068
rect 489236 31028 506480 31056
rect 489236 31016 489242 31028
rect 506474 31016 506480 31028
rect 506532 31016 506538 31068
rect 276106 29588 276112 29640
rect 276164 29628 276170 29640
rect 488534 29628 488540 29640
rect 276164 29600 488540 29628
rect 276164 29588 276170 29600
rect 488534 29588 488540 29600
rect 488592 29588 488598 29640
rect 143626 28228 143632 28280
rect 143684 28268 143690 28280
rect 353386 28268 353392 28280
rect 143684 28240 353392 28268
rect 143684 28228 143690 28240
rect 353386 28228 353392 28240
rect 353444 28228 353450 28280
rect 226426 25576 226432 25628
rect 226484 25616 226490 25628
rect 336734 25616 336740 25628
rect 226484 25588 336740 25616
rect 226484 25576 226490 25588
rect 336734 25576 336740 25588
rect 336792 25576 336798 25628
rect 230198 25508 230204 25560
rect 230256 25548 230262 25560
rect 343634 25548 343640 25560
rect 230256 25520 343640 25548
rect 230256 25508 230262 25520
rect 343634 25508 343640 25520
rect 343692 25508 343698 25560
rect 368474 25508 368480 25560
rect 368532 25548 368538 25560
rect 538214 25548 538220 25560
rect 368532 25520 538220 25548
rect 368532 25508 368538 25520
rect 538214 25508 538220 25520
rect 538272 25508 538278 25560
rect 161474 24080 161480 24132
rect 161532 24120 161538 24132
rect 379606 24120 379612 24132
rect 161532 24092 379612 24120
rect 161532 24080 161538 24092
rect 379606 24080 379612 24092
rect 379664 24080 379670 24132
rect 394786 24080 394792 24132
rect 394844 24120 394850 24132
rect 514754 24120 514760 24132
rect 394844 24092 514760 24120
rect 394844 24080 394850 24092
rect 514754 24080 514760 24092
rect 514812 24080 514818 24132
rect 3510 22720 3516 22772
rect 3568 22760 3574 22772
rect 189718 22760 189724 22772
rect 3568 22732 189724 22760
rect 3568 22720 3574 22732
rect 189718 22720 189724 22732
rect 189776 22720 189782 22772
rect 325694 22720 325700 22772
rect 325752 22760 325758 22772
rect 473446 22760 473452 22772
rect 325752 22732 473452 22760
rect 325752 22720 325758 22732
rect 473446 22720 473452 22732
rect 473504 22720 473510 22772
rect 168466 21360 168472 21412
rect 168524 21400 168530 21412
rect 307938 21400 307944 21412
rect 168524 21372 307944 21400
rect 168524 21360 168530 21372
rect 307938 21360 307944 21372
rect 307996 21360 308002 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 288434 20652 288440 20664
rect 3476 20624 288440 20652
rect 3476 20612 3482 20624
rect 288434 20612 288440 20624
rect 288492 20612 288498 20664
rect 538858 20612 538864 20664
rect 538916 20652 538922 20664
rect 579982 20652 579988 20664
rect 538916 20624 579988 20652
rect 538916 20612 538922 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 421006 18572 421012 18624
rect 421064 18612 421070 18624
rect 463970 18612 463976 18624
rect 421064 18584 463976 18612
rect 421064 18572 421070 18584
rect 463970 18572 463976 18584
rect 464028 18572 464034 18624
rect 367186 17212 367192 17264
rect 367244 17252 367250 17264
rect 392026 17252 392032 17264
rect 367244 17224 392032 17252
rect 367244 17212 367250 17224
rect 392026 17212 392032 17224
rect 392084 17212 392090 17264
rect 418246 17212 418252 17264
rect 418304 17252 418310 17264
rect 444466 17252 444472 17264
rect 418304 17224 444472 17252
rect 418304 17212 418310 17224
rect 444466 17212 444472 17224
rect 444524 17212 444530 17264
rect 371234 15852 371240 15904
rect 371292 15892 371298 15904
rect 533246 15892 533252 15904
rect 371292 15864 533252 15892
rect 371292 15852 371298 15864
rect 533246 15852 533252 15864
rect 533304 15852 533310 15904
rect 307846 14424 307852 14476
rect 307904 14464 307910 14476
rect 326338 14464 326344 14476
rect 307904 14436 326344 14464
rect 307904 14424 307910 14436
rect 326338 14424 326344 14436
rect 326396 14424 326402 14476
rect 465718 14424 465724 14476
rect 465776 14464 465782 14476
rect 509602 14464 509608 14476
rect 465776 14436 509608 14464
rect 465776 14424 465782 14436
rect 509602 14424 509608 14436
rect 509660 14424 509666 14476
rect 230382 13132 230388 13184
rect 230440 13172 230446 13184
rect 273346 13172 273352 13184
rect 230440 13144 273352 13172
rect 230440 13132 230446 13144
rect 273346 13132 273352 13144
rect 273404 13132 273410 13184
rect 110506 13064 110512 13116
rect 110564 13104 110570 13116
rect 167638 13104 167644 13116
rect 110564 13076 167644 13104
rect 110564 13064 110570 13076
rect 167638 13064 167644 13076
rect 167696 13064 167702 13116
rect 235810 13064 235816 13116
rect 235868 13104 235874 13116
rect 314654 13104 314660 13116
rect 235868 13076 314660 13104
rect 235868 13064 235874 13076
rect 314654 13064 314660 13076
rect 314712 13064 314718 13116
rect 357526 13064 357532 13116
rect 357584 13104 357590 13116
rect 544378 13104 544384 13116
rect 357584 13076 544384 13104
rect 357584 13064 357590 13076
rect 544378 13064 544384 13076
rect 544436 13064 544442 13116
rect 126974 11772 126980 11824
rect 127032 11812 127038 11824
rect 128170 11812 128176 11824
rect 127032 11784 128176 11812
rect 127032 11772 127038 11784
rect 128170 11772 128176 11784
rect 128228 11772 128234 11824
rect 184934 11772 184940 11824
rect 184992 11812 184998 11824
rect 186130 11812 186136 11824
rect 184992 11784 186136 11812
rect 184992 11772 184998 11784
rect 186130 11772 186136 11784
rect 186188 11772 186194 11824
rect 109034 11704 109040 11756
rect 109092 11744 109098 11756
rect 217318 11744 217324 11756
rect 109092 11716 217324 11744
rect 109092 11704 109098 11716
rect 217318 11704 217324 11716
rect 217376 11704 217382 11756
rect 227438 11704 227444 11756
rect 227496 11744 227502 11756
rect 227622 11744 227628 11756
rect 227496 11716 227628 11744
rect 227496 11704 227502 11716
rect 227622 11704 227628 11716
rect 227680 11704 227686 11756
rect 270586 11704 270592 11756
rect 270644 11744 270650 11756
rect 526162 11744 526168 11756
rect 270644 11716 526168 11744
rect 270644 11704 270650 11716
rect 526162 11704 526168 11716
rect 526220 11704 526226 11756
rect 77386 10276 77392 10328
rect 77444 10316 77450 10328
rect 220078 10316 220084 10328
rect 77444 10288 220084 10316
rect 77444 10276 77450 10288
rect 220078 10276 220084 10288
rect 220136 10276 220142 10328
rect 221090 10276 221096 10328
rect 221148 10316 221154 10328
rect 327074 10316 327080 10328
rect 221148 10288 327080 10316
rect 221148 10276 221154 10288
rect 327074 10276 327080 10288
rect 327132 10276 327138 10328
rect 331214 10276 331220 10328
rect 331272 10316 331278 10328
rect 515490 10316 515496 10328
rect 331272 10288 515496 10316
rect 331272 10276 331278 10288
rect 515490 10276 515496 10288
rect 515548 10276 515554 10328
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 464338 9596 464344 9648
rect 464396 9636 464402 9648
rect 465166 9636 465172 9648
rect 464396 9608 465172 9636
rect 464396 9596 464402 9608
rect 465166 9596 465172 9608
rect 465224 9596 465230 9648
rect 224862 9188 224868 9240
rect 224920 9228 224926 9240
rect 300762 9228 300768 9240
rect 224920 9200 300768 9228
rect 224920 9188 224926 9200
rect 300762 9188 300768 9200
rect 300820 9188 300826 9240
rect 228818 9120 228824 9172
rect 228876 9160 228882 9172
rect 362310 9160 362316 9172
rect 228876 9132 362316 9160
rect 228876 9120 228882 9132
rect 362310 9120 362316 9132
rect 362368 9120 362374 9172
rect 230290 9052 230296 9104
rect 230348 9092 230354 9104
rect 400122 9092 400128 9104
rect 230348 9064 400128 9092
rect 230348 9052 230354 9064
rect 400122 9052 400128 9064
rect 400180 9052 400186 9104
rect 73798 8984 73804 9036
rect 73856 9024 73862 9036
rect 224218 9024 224224 9036
rect 73856 8996 224224 9024
rect 73856 8984 73862 8996
rect 224218 8984 224224 8996
rect 224276 8984 224282 9036
rect 264974 8984 264980 9036
rect 265032 9024 265038 9036
rect 461670 9024 461676 9036
rect 265032 8996 461676 9024
rect 265032 8984 265038 8996
rect 461670 8984 461676 8996
rect 461728 8984 461734 9036
rect 222930 8916 222936 8968
rect 222988 8956 222994 8968
rect 426158 8956 426164 8968
rect 222988 8928 426164 8956
rect 222988 8916 222994 8928
rect 426158 8916 426164 8928
rect 426216 8916 426222 8968
rect 468478 8916 468484 8968
rect 468536 8956 468542 8968
rect 491110 8956 491116 8968
rect 468536 8928 491116 8956
rect 468536 8916 468542 8928
rect 491110 8916 491116 8928
rect 491168 8916 491174 8968
rect 502978 8916 502984 8968
rect 503036 8956 503042 8968
rect 520734 8956 520740 8968
rect 503036 8928 520740 8956
rect 503036 8916 503042 8928
rect 520734 8916 520740 8928
rect 520792 8916 520798 8968
rect 526438 8916 526444 8968
rect 526496 8956 526502 8968
rect 540790 8956 540796 8968
rect 526496 8928 540796 8956
rect 526496 8916 526502 8928
rect 540790 8916 540796 8928
rect 540848 8916 540854 8968
rect 273254 7964 273260 8016
rect 273312 8004 273318 8016
rect 301958 8004 301964 8016
rect 273312 7976 301964 8004
rect 273312 7964 273318 7976
rect 301958 7964 301964 7976
rect 302016 7964 302022 8016
rect 167178 7896 167184 7948
rect 167236 7936 167242 7948
rect 346394 7936 346400 7948
rect 167236 7908 346400 7936
rect 167236 7896 167242 7908
rect 346394 7896 346400 7908
rect 346452 7896 346458 7948
rect 112806 7828 112812 7880
rect 112864 7868 112870 7880
rect 304994 7868 305000 7880
rect 112864 7840 305000 7868
rect 112864 7828 112870 7840
rect 304994 7828 305000 7840
rect 305052 7828 305058 7880
rect 305546 7828 305552 7880
rect 305604 7868 305610 7880
rect 441706 7868 441712 7880
rect 305604 7840 441712 7868
rect 305604 7828 305610 7840
rect 441706 7828 441712 7840
rect 441764 7828 441770 7880
rect 291286 7760 291292 7812
rect 291344 7800 291350 7812
rect 507670 7800 507676 7812
rect 291344 7772 507676 7800
rect 291344 7760 291350 7772
rect 507670 7760 507676 7772
rect 507728 7760 507734 7812
rect 177850 7692 177856 7744
rect 177908 7732 177914 7744
rect 415486 7732 415492 7744
rect 177908 7704 415492 7732
rect 177908 7692 177914 7704
rect 415486 7692 415492 7704
rect 415544 7692 415550 7744
rect 277486 7624 277492 7676
rect 277544 7664 277550 7676
rect 543182 7664 543188 7676
rect 277544 7636 543188 7664
rect 277544 7624 277550 7636
rect 543182 7624 543188 7636
rect 543240 7624 543246 7676
rect 151906 7556 151912 7608
rect 151964 7596 151970 7608
rect 442994 7596 443000 7608
rect 151964 7568 443000 7596
rect 151964 7556 151970 7568
rect 442994 7556 443000 7568
rect 443052 7556 443058 7608
rect 549898 7556 549904 7608
rect 549956 7596 549962 7608
rect 562042 7596 562048 7608
rect 549956 7568 562048 7596
rect 549956 7556 549962 7568
rect 562042 7556 562048 7568
rect 562100 7556 562106 7608
rect 542998 6876 543004 6928
rect 543056 6916 543062 6928
rect 547874 6916 547880 6928
rect 543056 6888 547880 6916
rect 543056 6876 543062 6888
rect 547874 6876 547880 6888
rect 547932 6876 547938 6928
rect 222010 6808 222016 6860
rect 222068 6848 222074 6860
rect 306742 6848 306748 6860
rect 222068 6820 306748 6848
rect 222068 6808 222074 6820
rect 306742 6808 306748 6820
rect 306800 6808 306806 6860
rect 461578 6808 461584 6860
rect 461636 6848 461642 6860
rect 580166 6848 580172 6860
rect 461636 6820 580172 6848
rect 461636 6808 461642 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 227346 6740 227352 6792
rect 227404 6780 227410 6792
rect 313826 6780 313832 6792
rect 227404 6752 313832 6780
rect 227404 6740 227410 6752
rect 313826 6740 313832 6752
rect 313884 6740 313890 6792
rect 247586 6672 247592 6724
rect 247644 6712 247650 6724
rect 339494 6712 339500 6724
rect 247644 6684 339500 6712
rect 247644 6672 247650 6684
rect 339494 6672 339500 6684
rect 339552 6672 339558 6724
rect 206186 6604 206192 6656
rect 206244 6644 206250 6656
rect 299474 6644 299480 6656
rect 206244 6616 299480 6644
rect 206244 6604 206250 6616
rect 299474 6604 299480 6616
rect 299532 6604 299538 6656
rect 220722 6536 220728 6588
rect 220780 6576 220786 6588
rect 324406 6576 324412 6588
rect 220780 6548 324412 6576
rect 220780 6536 220786 6548
rect 324406 6536 324412 6548
rect 324464 6536 324470 6588
rect 354674 6536 354680 6588
rect 354732 6576 354738 6588
rect 385954 6576 385960 6588
rect 354732 6548 385960 6576
rect 354732 6536 354738 6548
rect 385954 6536 385960 6548
rect 386012 6536 386018 6588
rect 229830 6468 229836 6520
rect 229888 6508 229894 6520
rect 335354 6508 335360 6520
rect 229888 6480 335360 6508
rect 229888 6468 229894 6480
rect 335354 6468 335360 6480
rect 335412 6468 335418 6520
rect 357526 6468 357532 6520
rect 357584 6508 357590 6520
rect 408494 6508 408500 6520
rect 357584 6480 408500 6508
rect 357584 6468 357590 6480
rect 408494 6468 408500 6480
rect 408552 6468 408558 6520
rect 216582 6400 216588 6452
rect 216640 6440 216646 6452
rect 363506 6440 363512 6452
rect 216640 6412 363512 6440
rect 216640 6400 216646 6412
rect 363506 6400 363512 6412
rect 363564 6400 363570 6452
rect 375282 6400 375288 6452
rect 375340 6440 375346 6452
rect 391934 6440 391940 6452
rect 375340 6412 391940 6440
rect 375340 6400 375346 6412
rect 391934 6400 391940 6412
rect 391992 6400 391998 6452
rect 131758 6332 131764 6384
rect 131816 6372 131822 6384
rect 296806 6372 296812 6384
rect 131816 6344 296812 6372
rect 131816 6332 131822 6344
rect 296806 6332 296812 6344
rect 296864 6332 296870 6384
rect 302326 6332 302332 6384
rect 302384 6372 302390 6384
rect 322106 6372 322112 6384
rect 302384 6344 322112 6372
rect 302384 6332 302390 6344
rect 322106 6332 322112 6344
rect 322164 6332 322170 6384
rect 361114 6332 361120 6384
rect 361172 6372 361178 6384
rect 429286 6372 429292 6384
rect 361172 6344 429292 6372
rect 361172 6332 361178 6344
rect 429286 6332 429292 6344
rect 429344 6332 429350 6384
rect 220538 6264 220544 6316
rect 220596 6304 220602 6316
rect 255866 6304 255872 6316
rect 220596 6276 255872 6304
rect 220596 6264 220602 6276
rect 255866 6264 255872 6276
rect 255924 6264 255930 6316
rect 258258 6264 258264 6316
rect 258316 6304 258322 6316
rect 430666 6304 430672 6316
rect 258316 6276 430672 6304
rect 258316 6264 258322 6276
rect 430666 6264 430672 6276
rect 430724 6264 430730 6316
rect 224494 6196 224500 6248
rect 224552 6236 224558 6248
rect 407206 6236 407212 6248
rect 224552 6208 407212 6236
rect 224552 6196 224558 6208
rect 407206 6196 407212 6208
rect 407264 6196 407270 6248
rect 134150 6128 134156 6180
rect 134208 6168 134214 6180
rect 393314 6168 393320 6180
rect 134208 6140 393320 6168
rect 134208 6128 134214 6140
rect 393314 6128 393320 6140
rect 393372 6128 393378 6180
rect 220630 6060 220636 6112
rect 220688 6100 220694 6112
rect 296070 6100 296076 6112
rect 220688 6072 296076 6100
rect 220688 6060 220694 6072
rect 296070 6060 296076 6072
rect 296128 6060 296134 6112
rect 223482 5992 223488 6044
rect 223540 6032 223546 6044
rect 276014 6032 276020 6044
rect 223540 6004 276020 6032
rect 223540 5992 223546 6004
rect 276014 5992 276020 6004
rect 276072 5992 276078 6044
rect 223022 5924 223028 5976
rect 223080 5964 223086 5976
rect 252370 5964 252376 5976
rect 223080 5936 252376 5964
rect 223080 5924 223086 5936
rect 252370 5924 252376 5936
rect 252428 5924 252434 5976
rect 256694 5924 256700 5976
rect 256752 5964 256758 5976
rect 293678 5964 293684 5976
rect 256752 5936 293684 5964
rect 256752 5924 256758 5936
rect 293678 5924 293684 5936
rect 293736 5924 293742 5976
rect 436738 5516 436744 5568
rect 436796 5556 436802 5568
rect 443822 5556 443828 5568
rect 436796 5528 443828 5556
rect 436796 5516 436802 5528
rect 443822 5516 443828 5528
rect 443880 5516 443886 5568
rect 227438 5380 227444 5432
rect 227496 5420 227502 5432
rect 227622 5420 227628 5432
rect 227496 5392 227628 5420
rect 227496 5380 227502 5392
rect 227622 5380 227628 5392
rect 227680 5380 227686 5432
rect 339862 5176 339868 5228
rect 339920 5216 339926 5228
rect 350534 5216 350540 5228
rect 339920 5188 350540 5216
rect 339920 5176 339926 5188
rect 350534 5176 350540 5188
rect 350592 5176 350598 5228
rect 238846 5108 238852 5160
rect 238904 5148 238910 5160
rect 274818 5148 274824 5160
rect 238904 5120 274824 5148
rect 238904 5108 238910 5120
rect 274818 5108 274824 5120
rect 274876 5108 274882 5160
rect 307938 5108 307944 5160
rect 307996 5148 308002 5160
rect 356054 5148 356060 5160
rect 307996 5120 356060 5148
rect 307996 5108 308002 5120
rect 356054 5108 356060 5120
rect 356112 5108 356118 5160
rect 220446 5040 220452 5092
rect 220504 5080 220510 5092
rect 258074 5080 258080 5092
rect 220504 5052 258080 5080
rect 220504 5040 220510 5052
rect 258074 5040 258080 5052
rect 258132 5040 258138 5092
rect 286594 5040 286600 5092
rect 286652 5080 286658 5092
rect 358906 5080 358912 5092
rect 286652 5052 358912 5080
rect 286652 5040 286658 5052
rect 358906 5040 358912 5052
rect 358964 5040 358970 5092
rect 202690 4972 202696 5024
rect 202748 5012 202754 5024
rect 248506 5012 248512 5024
rect 202748 4984 248512 5012
rect 202748 4972 202754 4984
rect 248506 4972 248512 4984
rect 248564 4972 248570 5024
rect 257062 4972 257068 5024
rect 257120 5012 257126 5024
rect 332594 5012 332600 5024
rect 257120 4984 332600 5012
rect 257120 4972 257126 4984
rect 332594 4972 332600 4984
rect 332652 4972 332658 5024
rect 347866 4972 347872 5024
rect 347924 5012 347930 5024
rect 402514 5012 402520 5024
rect 347924 4984 402520 5012
rect 347924 4972 347930 4984
rect 402514 4972 402520 4984
rect 402572 4972 402578 5024
rect 236086 4904 236092 4956
rect 236144 4944 236150 4956
rect 317322 4944 317328 4956
rect 236144 4916 317328 4944
rect 236144 4904 236150 4916
rect 317322 4904 317328 4916
rect 317380 4904 317386 4956
rect 338666 4904 338672 4956
rect 338724 4944 338730 4956
rect 409966 4944 409972 4956
rect 338724 4916 409972 4944
rect 338724 4904 338730 4916
rect 409966 4904 409972 4916
rect 410024 4904 410030 4956
rect 53742 4836 53748 4888
rect 53800 4876 53806 4888
rect 240226 4876 240232 4888
rect 53800 4848 240232 4876
rect 53800 4836 53806 4848
rect 240226 4836 240232 4848
rect 240284 4836 240290 4888
rect 253474 4836 253480 4888
rect 253532 4876 253538 4888
rect 407298 4876 407304 4888
rect 253532 4848 407304 4876
rect 253532 4836 253538 4848
rect 407298 4836 407304 4848
rect 407356 4836 407362 4888
rect 414014 4836 414020 4888
rect 414072 4876 414078 4888
rect 432046 4876 432052 4888
rect 414072 4848 432052 4876
rect 414072 4836 414078 4848
rect 432046 4836 432052 4848
rect 432104 4836 432110 4888
rect 140038 4768 140044 4820
rect 140096 4808 140102 4820
rect 372614 4808 372620 4820
rect 140096 4780 372620 4808
rect 140096 4768 140102 4780
rect 372614 4768 372620 4780
rect 372672 4768 372678 4820
rect 413094 4768 413100 4820
rect 413152 4808 413158 4820
rect 444374 4808 444380 4820
rect 413152 4780 444380 4808
rect 413152 4768 413158 4780
rect 444374 4768 444380 4780
rect 444432 4768 444438 4820
rect 476758 4768 476764 4820
rect 476816 4808 476822 4820
rect 499390 4808 499396 4820
rect 476816 4780 499396 4808
rect 476816 4768 476822 4780
rect 499390 4768 499396 4780
rect 499448 4768 499454 4820
rect 227456 4168 227760 4196
rect 223390 4020 223396 4072
rect 223448 4060 223454 4072
rect 227456 4060 227484 4168
rect 227732 4128 227760 4168
rect 422294 4156 422300 4208
rect 422352 4196 422358 4208
rect 423766 4196 423772 4208
rect 422352 4168 423772 4196
rect 422352 4156 422358 4168
rect 423766 4156 423772 4168
rect 423824 4156 423830 4208
rect 544470 4156 544476 4208
rect 544528 4196 544534 4208
rect 545482 4196 545488 4208
rect 544528 4168 545488 4196
rect 544528 4156 544534 4168
rect 545482 4156 545488 4168
rect 545540 4156 545546 4208
rect 264146 4128 264152 4140
rect 227732 4100 264152 4128
rect 264146 4088 264152 4100
rect 264204 4088 264210 4140
rect 434438 4088 434444 4140
rect 434496 4128 434502 4140
rect 462406 4128 462412 4140
rect 434496 4100 462412 4128
rect 434496 4088 434502 4100
rect 462406 4088 462412 4100
rect 462464 4088 462470 4140
rect 475378 4088 475384 4140
rect 475436 4128 475442 4140
rect 475930 4128 475936 4140
rect 475436 4100 475936 4128
rect 475436 4088 475442 4100
rect 475930 4088 475936 4100
rect 475988 4088 475994 4140
rect 223448 4032 227484 4060
rect 223448 4020 223454 4032
rect 227530 4020 227536 4072
rect 227588 4060 227594 4072
rect 288986 4060 288992 4072
rect 227588 4032 288992 4060
rect 227588 4020 227594 4032
rect 288986 4020 288992 4032
rect 289044 4020 289050 4072
rect 427262 4020 427268 4072
rect 427320 4060 427326 4072
rect 459554 4060 459560 4072
rect 427320 4032 459560 4060
rect 427320 4020 427326 4032
rect 459554 4020 459560 4032
rect 459612 4020 459618 4072
rect 227254 3952 227260 4004
rect 227312 3992 227318 4004
rect 290182 3992 290188 4004
rect 227312 3964 290188 3992
rect 227312 3952 227318 3964
rect 290182 3952 290188 3964
rect 290240 3952 290246 4004
rect 414290 3952 414296 4004
rect 414348 3992 414354 4004
rect 461026 3992 461032 4004
rect 414348 3964 461032 3992
rect 414348 3952 414354 3964
rect 461026 3952 461032 3964
rect 461084 3952 461090 4004
rect 225414 3884 225420 3936
rect 225472 3924 225478 3936
rect 227346 3924 227352 3936
rect 225472 3896 227352 3924
rect 225472 3884 225478 3896
rect 227346 3884 227352 3896
rect 227404 3884 227410 3936
rect 227714 3884 227720 3936
rect 227772 3924 227778 3936
rect 299658 3924 299664 3936
rect 227772 3896 299664 3924
rect 227772 3884 227778 3896
rect 299658 3884 299664 3896
rect 299716 3884 299722 3936
rect 416682 3884 416688 3936
rect 416740 3924 416746 3936
rect 463878 3924 463884 3936
rect 416740 3896 463884 3924
rect 416740 3884 416746 3896
rect 463878 3884 463884 3896
rect 463936 3884 463942 3936
rect 226150 3816 226156 3868
rect 226208 3856 226214 3868
rect 332594 3856 332600 3868
rect 226208 3828 332600 3856
rect 226208 3816 226214 3828
rect 332594 3816 332600 3828
rect 332652 3816 332658 3868
rect 367830 3816 367836 3868
rect 367888 3856 367894 3868
rect 459186 3856 459192 3868
rect 367888 3828 459192 3856
rect 367888 3816 367894 3828
rect 459186 3816 459192 3828
rect 459244 3816 459250 3868
rect 135254 3748 135260 3800
rect 135312 3788 135318 3800
rect 136450 3788 136456 3800
rect 135312 3760 136456 3788
rect 135312 3748 135318 3760
rect 136450 3748 136456 3760
rect 136508 3748 136514 3800
rect 151814 3748 151820 3800
rect 151872 3788 151878 3800
rect 153010 3788 153016 3800
rect 151872 3760 153016 3788
rect 151872 3748 151878 3760
rect 153010 3748 153016 3760
rect 153068 3748 153074 3800
rect 193214 3748 193220 3800
rect 193272 3788 193278 3800
rect 194410 3788 194416 3800
rect 193272 3760 194416 3788
rect 193272 3748 193278 3760
rect 194410 3748 194416 3760
rect 194468 3748 194474 3800
rect 226334 3748 226340 3800
rect 226392 3788 226398 3800
rect 227530 3788 227536 3800
rect 226392 3760 227536 3788
rect 226392 3748 226398 3760
rect 227530 3748 227536 3760
rect 227588 3748 227594 3800
rect 227622 3748 227628 3800
rect 227680 3788 227686 3800
rect 371694 3788 371700 3800
rect 227680 3760 371700 3788
rect 227680 3748 227686 3760
rect 371694 3748 371700 3760
rect 371752 3748 371758 3800
rect 404814 3748 404820 3800
rect 404872 3788 404878 3800
rect 459738 3788 459744 3800
rect 404872 3760 459744 3788
rect 404872 3748 404878 3760
rect 459738 3748 459744 3760
rect 459796 3748 459802 3800
rect 525058 3748 525064 3800
rect 525116 3788 525122 3800
rect 557350 3788 557356 3800
rect 525116 3760 557356 3788
rect 525116 3748 525122 3760
rect 557350 3748 557356 3760
rect 557408 3748 557414 3800
rect 103330 3680 103336 3732
rect 103388 3720 103394 3732
rect 249886 3720 249892 3732
rect 103388 3692 249892 3720
rect 103388 3680 103394 3692
rect 249886 3680 249892 3692
rect 249944 3680 249950 3732
rect 265342 3680 265348 3732
rect 265400 3720 265406 3732
rect 450538 3720 450544 3732
rect 265400 3692 450544 3720
rect 265400 3680 265406 3692
rect 450538 3680 450544 3692
rect 450596 3680 450602 3732
rect 455690 3680 455696 3732
rect 455748 3720 455754 3732
rect 462590 3720 462596 3732
rect 455748 3692 462596 3720
rect 455748 3680 455754 3692
rect 462590 3680 462596 3692
rect 462648 3680 462654 3732
rect 500218 3680 500224 3732
rect 500276 3720 500282 3732
rect 532510 3720 532516 3732
rect 500276 3692 532516 3720
rect 500276 3680 500282 3692
rect 532510 3680 532516 3692
rect 532568 3680 532574 3732
rect 533338 3680 533344 3732
rect 533396 3720 533402 3732
rect 536098 3720 536104 3732
rect 533396 3692 536104 3720
rect 533396 3680 533402 3692
rect 536098 3680 536104 3692
rect 536156 3680 536162 3732
rect 114002 3612 114008 3664
rect 114060 3652 114066 3664
rect 351914 3652 351920 3664
rect 114060 3624 351920 3652
rect 114060 3612 114066 3624
rect 351914 3612 351920 3624
rect 351972 3612 351978 3664
rect 355226 3612 355232 3664
rect 355284 3652 355290 3664
rect 460934 3652 460940 3664
rect 355284 3624 460940 3652
rect 355284 3612 355290 3624
rect 460934 3612 460940 3624
rect 460992 3612 460998 3664
rect 504358 3612 504364 3664
rect 504416 3652 504422 3664
rect 539594 3652 539600 3664
rect 504416 3624 539600 3652
rect 504416 3612 504422 3624
rect 539594 3612 539600 3624
rect 539652 3612 539658 3664
rect 555418 3612 555424 3664
rect 555476 3652 555482 3664
rect 565630 3652 565636 3664
rect 555476 3624 565636 3652
rect 555476 3612 555482 3624
rect 565630 3612 565636 3624
rect 565688 3612 565694 3664
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 280798 3584 280804 3596
rect 24268 3556 280804 3584
rect 24268 3544 24274 3556
rect 280798 3544 280804 3556
rect 280856 3544 280862 3596
rect 315022 3544 315028 3596
rect 315080 3584 315086 3596
rect 446398 3584 446404 3596
rect 315080 3556 446404 3584
rect 315080 3544 315086 3556
rect 446398 3544 446404 3556
rect 446456 3544 446462 3596
rect 447778 3544 447784 3596
rect 447836 3584 447842 3596
rect 448606 3584 448612 3596
rect 447836 3556 448612 3584
rect 447836 3544 447842 3556
rect 448606 3544 448612 3556
rect 448664 3544 448670 3596
rect 453298 3544 453304 3596
rect 453356 3584 453362 3596
rect 461118 3584 461124 3596
rect 453356 3556 461124 3584
rect 453356 3544 453362 3556
rect 461118 3544 461124 3556
rect 461176 3544 461182 3596
rect 471238 3544 471244 3596
rect 471296 3584 471302 3596
rect 486418 3584 486424 3596
rect 471296 3556 486424 3584
rect 471296 3544 471302 3556
rect 486418 3544 486424 3556
rect 486476 3544 486482 3596
rect 486510 3544 486516 3596
rect 486568 3584 486574 3596
rect 500586 3584 500592 3596
rect 486568 3556 500592 3584
rect 486568 3544 486574 3556
rect 500586 3544 500592 3556
rect 500644 3544 500650 3596
rect 520918 3544 520924 3596
rect 520976 3584 520982 3596
rect 563238 3584 563244 3596
rect 520976 3556 563244 3584
rect 520976 3544 520982 3556
rect 563238 3544 563244 3556
rect 563296 3544 563302 3596
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3694 3516 3700 3528
rect 2832 3488 3700 3516
rect 2832 3476 2838 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11980 3516
rect 11112 3476 11118 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 21358 3516 21364 3528
rect 13596 3488 21364 3516
rect 13596 3476 13602 3488
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 28902 3476 28908 3528
rect 28960 3516 28966 3528
rect 317414 3516 317420 3528
rect 28960 3488 317420 3516
rect 28960 3476 28966 3488
rect 317414 3476 317420 3488
rect 317472 3476 317478 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 332686 3476 332692 3528
rect 332744 3516 332750 3528
rect 333882 3516 333888 3528
rect 332744 3488 333888 3516
rect 332744 3476 332750 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 340874 3476 340880 3528
rect 340932 3516 340938 3528
rect 342162 3516 342168 3528
rect 340932 3488 342168 3516
rect 340932 3476 340938 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 350442 3476 350448 3528
rect 350500 3516 350506 3528
rect 453574 3516 453580 3528
rect 350500 3488 453580 3516
rect 350500 3476 350506 3488
rect 453574 3476 453580 3488
rect 453632 3476 453638 3528
rect 456886 3476 456892 3528
rect 456944 3516 456950 3528
rect 458082 3516 458088 3528
rect 456944 3488 458088 3516
rect 456944 3476 456950 3488
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 460198 3476 460204 3528
rect 460256 3516 460262 3528
rect 546678 3516 546684 3528
rect 460256 3488 546684 3516
rect 460256 3476 460262 3488
rect 546678 3476 546684 3488
rect 546736 3476 546742 3528
rect 562318 3476 562324 3528
rect 562376 3516 562382 3528
rect 576302 3516 576308 3528
rect 562376 3488 576308 3516
rect 562376 3476 562382 3488
rect 576302 3476 576308 3488
rect 576360 3476 576366 3528
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 26878 3448 26884 3460
rect 18288 3420 26884 3448
rect 18288 3408 18294 3420
rect 26878 3408 26884 3420
rect 26936 3408 26942 3460
rect 44174 3408 44180 3460
rect 44232 3448 44238 3460
rect 45094 3448 45100 3460
rect 44232 3420 45100 3448
rect 44232 3408 44238 3420
rect 45094 3408 45100 3420
rect 45152 3408 45158 3460
rect 69014 3408 69020 3460
rect 69072 3448 69078 3460
rect 69934 3448 69940 3460
rect 69072 3420 69940 3448
rect 69072 3408 69078 3420
rect 69934 3408 69940 3420
rect 69992 3408 69998 3460
rect 77294 3408 77300 3460
rect 77352 3448 77358 3460
rect 78214 3448 78220 3460
rect 77352 3420 78220 3448
rect 77352 3408 77358 3420
rect 78214 3408 78220 3420
rect 78272 3408 78278 3460
rect 93854 3408 93860 3460
rect 93912 3448 93918 3460
rect 94774 3448 94780 3460
rect 93912 3420 94780 3448
rect 93912 3408 93918 3420
rect 94774 3408 94780 3420
rect 94832 3408 94838 3460
rect 110414 3408 110420 3460
rect 110472 3448 110478 3460
rect 111610 3448 111616 3460
rect 110472 3420 111616 3448
rect 110472 3408 110478 3420
rect 111610 3408 111616 3420
rect 111668 3408 111674 3460
rect 161290 3408 161296 3460
rect 161348 3448 161354 3460
rect 226978 3448 226984 3460
rect 161348 3420 226984 3448
rect 161348 3408 161354 3420
rect 226978 3408 226984 3420
rect 227036 3408 227042 3460
rect 228358 3408 228364 3460
rect 228416 3448 228422 3460
rect 523034 3448 523040 3460
rect 228416 3420 523040 3448
rect 228416 3408 228422 3420
rect 523034 3408 523040 3420
rect 523092 3408 523098 3460
rect 529198 3408 529204 3460
rect 529256 3448 529262 3460
rect 564434 3448 564440 3460
rect 529256 3420 564440 3448
rect 529256 3408 529262 3420
rect 564434 3408 564440 3420
rect 564492 3408 564498 3460
rect 21818 3340 21824 3392
rect 21876 3380 21882 3392
rect 28258 3380 28264 3392
rect 21876 3352 28264 3380
rect 21876 3340 21882 3352
rect 28258 3340 28264 3352
rect 28316 3340 28322 3392
rect 226058 3340 226064 3392
rect 226116 3380 226122 3392
rect 260650 3380 260656 3392
rect 226116 3352 260656 3380
rect 226116 3340 226122 3352
rect 260650 3340 260656 3352
rect 260708 3340 260714 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 367002 3380 367008 3392
rect 365772 3352 367008 3380
rect 365772 3340 365778 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 407114 3340 407120 3392
rect 407172 3380 407178 3392
rect 408402 3380 408408 3392
rect 407172 3352 408408 3380
rect 407172 3340 407178 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 423674 3340 423680 3392
rect 423732 3380 423738 3392
rect 424962 3380 424968 3392
rect 423732 3352 424968 3380
rect 423732 3340 423738 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 441522 3340 441528 3392
rect 441580 3380 441586 3392
rect 462498 3380 462504 3392
rect 441580 3352 462504 3380
rect 441580 3340 441586 3352
rect 462498 3340 462504 3352
rect 462556 3340 462562 3392
rect 576118 3340 576124 3392
rect 576176 3380 576182 3392
rect 577406 3380 577412 3392
rect 576176 3352 577412 3380
rect 576176 3340 576182 3352
rect 577406 3340 577412 3352
rect 577464 3340 577470 3392
rect 222102 3272 222108 3324
rect 222160 3312 222166 3324
rect 246390 3312 246396 3324
rect 222160 3284 246396 3312
rect 222160 3272 222166 3284
rect 246390 3272 246396 3284
rect 246448 3272 246454 3324
rect 446398 3272 446404 3324
rect 446456 3312 446462 3324
rect 452378 3312 452384 3324
rect 446456 3284 452384 3312
rect 446456 3272 446462 3284
rect 452378 3272 452384 3284
rect 452436 3272 452442 3324
rect 453574 3272 453580 3324
rect 453632 3312 453638 3324
rect 459002 3312 459008 3324
rect 453632 3284 459008 3312
rect 453632 3272 453638 3284
rect 459002 3272 459008 3284
rect 459060 3272 459066 3324
rect 475930 3272 475936 3324
rect 475988 3312 475994 3324
rect 481726 3312 481732 3324
rect 475988 3284 481732 3312
rect 475988 3272 475994 3284
rect 481726 3272 481732 3284
rect 481784 3272 481790 3324
rect 567838 3272 567844 3324
rect 567896 3312 567902 3324
rect 571518 3312 571524 3324
rect 567896 3284 571524 3312
rect 567896 3272 567902 3284
rect 571518 3272 571524 3284
rect 571576 3272 571582 3324
rect 571978 3272 571984 3324
rect 572036 3312 572042 3324
rect 572714 3312 572720 3324
rect 572036 3284 572720 3312
rect 572036 3272 572042 3284
rect 572714 3272 572720 3284
rect 572772 3272 572778 3324
rect 223206 3204 223212 3256
rect 223264 3244 223270 3256
rect 242894 3244 242900 3256
rect 223264 3216 242900 3244
rect 223264 3204 223270 3216
rect 242894 3204 242900 3216
rect 242952 3204 242958 3256
rect 449802 3204 449808 3256
rect 449860 3244 449866 3256
rect 465074 3244 465080 3256
rect 449860 3216 465080 3244
rect 449860 3204 449866 3216
rect 465074 3204 465080 3216
rect 465132 3204 465138 3256
rect 222746 3136 222752 3188
rect 222804 3176 222810 3188
rect 225598 3176 225604 3188
rect 222804 3148 225604 3176
rect 222804 3136 222810 3148
rect 225598 3136 225604 3148
rect 225656 3136 225662 3188
rect 450906 3136 450912 3188
rect 450964 3176 450970 3188
rect 464522 3176 464528 3188
rect 450964 3148 464528 3176
rect 450964 3136 450970 3148
rect 464522 3136 464528 3148
rect 464580 3136 464586 3188
rect 17034 3068 17040 3120
rect 17092 3108 17098 3120
rect 24118 3108 24124 3120
rect 17092 3080 24124 3108
rect 17092 3068 17098 3080
rect 24118 3068 24124 3080
rect 24176 3068 24182 3120
rect 433242 3068 433248 3120
rect 433300 3108 433306 3120
rect 451918 3108 451924 3120
rect 433300 3080 451924 3108
rect 433300 3068 433306 3080
rect 451918 3068 451924 3080
rect 451976 3068 451982 3120
rect 472618 3000 472624 3052
rect 472676 3040 472682 3052
rect 474550 3040 474556 3052
rect 472676 3012 474556 3040
rect 472676 3000 472682 3012
rect 474550 3000 474556 3012
rect 474608 3000 474614 3052
rect 548518 3000 548524 3052
rect 548576 3040 548582 3052
rect 554958 3040 554964 3052
rect 548576 3012 554964 3040
rect 548576 3000 548582 3012
rect 554958 3000 554964 3012
rect 555016 3000 555022 3052
rect 307754 2864 307760 2916
rect 307812 2904 307818 2916
rect 309042 2904 309048 2916
rect 307812 2876 309048 2904
rect 307812 2864 307818 2876
rect 309042 2864 309048 2876
rect 309100 2864 309106 2916
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 397460 700476 397512 700528
rect 459652 700476 459704 700528
rect 137836 700408 137888 700460
rect 157984 700408 158036 700460
rect 255320 700408 255372 700460
rect 332508 700408 332560 700460
rect 407120 700408 407172 700460
rect 543464 700408 543516 700460
rect 8116 700340 8168 700392
rect 131764 700340 131816 700392
rect 154120 700340 154172 700392
rect 256700 700340 256752 700392
rect 267648 700340 267700 700392
rect 436100 700340 436152 700392
rect 89168 700272 89220 700324
rect 227076 700272 227128 700324
rect 233976 700272 234028 700324
rect 527180 700272 527232 700324
rect 300124 699660 300176 699712
rect 306380 699660 306432 699712
rect 461676 699660 461728 699712
rect 462320 699660 462372 699712
rect 465724 696940 465776 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 340880 683136 340932 683188
rect 498844 683136 498896 683188
rect 580172 683136 580224 683188
rect 298100 670760 298152 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 452660 670692 452712 670744
rect 3424 656888 3476 656940
rect 79324 656888 79376 656940
rect 502984 643084 503036 643136
rect 580172 643084 580224 643136
rect 237380 630640 237432 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 314660 618264 314712 618316
rect 293960 616836 294012 616888
rect 580172 616836 580224 616888
rect 485044 590656 485096 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 21364 579640 21416 579692
rect 3424 577464 3476 577516
rect 453120 577464 453172 577516
rect 305460 574744 305512 574796
rect 429200 574744 429252 574796
rect 234252 571956 234304 572008
rect 412640 571956 412692 572008
rect 282920 570664 282972 570716
rect 453028 570664 453080 570716
rect 234160 570596 234212 570648
rect 580356 570596 580408 570648
rect 169760 566448 169812 566500
rect 453212 566448 453264 566500
rect 3424 565836 3476 565888
rect 345388 565836 345440 565888
rect 234344 563728 234396 563780
rect 347780 563728 347832 563780
rect 233148 563660 233200 563712
rect 364340 563660 364392 563712
rect 406568 563048 406620 563100
rect 579804 563048 579856 563100
rect 224316 562504 224368 562556
rect 371792 562504 371844 562556
rect 215300 562436 215352 562488
rect 426532 562436 426584 562488
rect 234528 562368 234580 562420
rect 494060 562368 494112 562420
rect 104900 562300 104952 562352
rect 456984 562300 457036 562352
rect 220452 562232 220504 562284
rect 441620 562232 441672 562284
rect 106280 562164 106332 562216
rect 340236 562164 340288 562216
rect 238760 562096 238812 562148
rect 500960 562096 501012 562148
rect 253296 562028 253348 562080
rect 531412 562028 531464 562080
rect 260380 561960 260432 562012
rect 540980 561960 541032 562012
rect 279056 561892 279108 561944
rect 572812 561892 572864 561944
rect 225972 561824 226024 561876
rect 270684 561824 270736 561876
rect 273260 561824 273312 561876
rect 576124 561824 576176 561876
rect 6920 561756 6972 561808
rect 324320 561756 324372 561808
rect 241704 561688 241756 561740
rect 569960 561688 570012 561740
rect 222844 561008 222896 561060
rect 350540 561008 350592 561060
rect 252008 560940 252060 560992
rect 558920 560940 558972 560992
rect 200764 560872 200816 560924
rect 316040 560872 316092 560924
rect 329288 560872 329340 560924
rect 483020 560872 483072 560924
rect 309324 560804 309376 560856
rect 465816 560804 465868 560856
rect 227352 560736 227404 560788
rect 271972 560736 272024 560788
rect 293224 560736 293276 560788
rect 464528 560736 464580 560788
rect 206284 560668 206336 560720
rect 382740 560668 382792 560720
rect 220176 560600 220228 560652
rect 268108 560600 268160 560652
rect 302884 560600 302936 560652
rect 480260 560600 480312 560652
rect 199384 560532 199436 560584
rect 280344 560532 280396 560584
rect 300308 560532 300360 560584
rect 487160 560532 487212 560584
rect 334440 560464 334492 560516
rect 538864 560464 538916 560516
rect 244280 560396 244332 560448
rect 507124 560396 507176 560448
rect 249800 560328 249852 560380
rect 527824 560328 527876 560380
rect 8944 560260 8996 560312
rect 445208 560260 445260 560312
rect 360936 559920 360988 559972
rect 446588 559920 446640 559972
rect 234896 559852 234948 559904
rect 368020 559852 368072 559904
rect 388628 559852 388680 559904
rect 451740 559852 451792 559904
rect 232412 559784 232464 559836
rect 393412 559784 393464 559836
rect 234712 559716 234764 559768
rect 424048 559716 424100 559768
rect 223488 559648 223540 559700
rect 245660 559648 245712 559700
rect 261668 559648 261720 559700
rect 301688 559648 301740 559700
rect 419448 559648 419500 559700
rect 459928 559648 459980 559700
rect 228364 559580 228416 559632
rect 289452 559580 289504 559632
rect 416688 559580 416740 559632
rect 461400 559580 461452 559632
rect 226800 559512 226852 559564
rect 288440 559512 288492 559564
rect 414388 559512 414440 559564
rect 460940 559512 460992 559564
rect 217324 559444 217376 559496
rect 263048 559444 263100 559496
rect 274732 559444 274784 559496
rect 362960 559444 363012 559496
rect 412456 559444 412508 559496
rect 459008 559444 459060 559496
rect 229928 559376 229980 559428
rect 322940 559376 322992 559428
rect 420828 559376 420880 559428
rect 457076 559376 457128 559428
rect 167644 559308 167696 559360
rect 292028 559308 292080 559360
rect 402152 559308 402204 559360
rect 456892 559308 456944 559360
rect 224224 559240 224276 559292
rect 354680 559240 354732 559292
rect 438216 559240 438268 559292
rect 465356 559240 465408 559292
rect 367008 559172 367060 559224
rect 389272 559172 389324 559224
rect 403440 559172 403492 559224
rect 458364 559172 458416 559224
rect 235816 559104 235868 559156
rect 378968 559104 379020 559156
rect 392492 559104 392544 559156
rect 451648 559104 451700 559156
rect 228456 559036 228508 559088
rect 377680 559036 377732 559088
rect 378784 559036 378836 559088
rect 430580 559036 430632 559088
rect 432420 559036 432472 559088
rect 464068 559036 464120 559088
rect 235908 558968 235960 559020
rect 261760 558968 261812 559020
rect 262864 558968 262916 559020
rect 274640 558968 274692 559020
rect 398288 558968 398340 559020
rect 462412 558968 462464 559020
rect 232780 558900 232832 558952
rect 265624 558900 265676 558952
rect 393320 558900 393372 558952
rect 421472 558900 421524 558952
rect 423404 558900 423456 558952
rect 469864 558900 469916 558952
rect 225604 558424 225656 558476
rect 284300 558424 284352 558476
rect 225420 558356 225472 558408
rect 287060 558356 287112 558408
rect 155960 558288 156012 558340
rect 274732 558288 274784 558340
rect 46940 558220 46992 558272
rect 262864 558220 262916 558272
rect 343548 558220 343600 558272
rect 453304 558220 453356 558272
rect 3424 558152 3476 558204
rect 378784 558152 378836 558204
rect 400864 558152 400916 558204
rect 481732 558152 481784 558204
rect 233884 558084 233936 558136
rect 320364 558084 320416 558136
rect 349988 558084 350040 558136
rect 460204 558084 460256 558136
rect 232872 558016 232924 558068
rect 328092 558016 328144 558068
rect 449808 558016 449860 558068
rect 472624 558016 472676 558068
rect 187700 557948 187752 558000
rect 356428 557948 356480 558000
rect 404728 557948 404780 558000
rect 503720 557948 503772 558000
rect 136640 557880 136692 557932
rect 317788 557880 317840 557932
rect 344836 557880 344888 557932
rect 466460 557880 466512 557932
rect 92480 557812 92532 557864
rect 285680 557812 285732 557864
rect 391204 557812 391256 557864
rect 524420 557812 524472 557864
rect 15200 557744 15252 557796
rect 259460 557744 259512 557796
rect 308772 557744 308824 557796
rect 465172 557744 465224 557796
rect 241152 557676 241204 557728
rect 492680 557676 492732 557728
rect 162860 557608 162912 557660
rect 433708 557608 433760 557660
rect 443368 557608 443420 557660
rect 496820 557608 496872 557660
rect 126980 557540 127032 557592
rect 405372 557540 405424 557592
rect 435640 557540 435692 557592
rect 565820 557540 565872 557592
rect 197360 557132 197412 557184
rect 353300 557132 353352 557184
rect 143540 557064 143592 557116
rect 369308 557064 369360 557116
rect 386052 557064 386104 557116
rect 453580 557064 453632 557116
rect 127072 556996 127124 557048
rect 366732 556996 366784 557048
rect 376668 556996 376720 557048
rect 451556 556996 451608 557048
rect 226156 556928 226208 556980
rect 266912 556928 266964 556980
rect 387340 556928 387392 556980
rect 469220 556928 469272 556980
rect 175280 556860 175332 556912
rect 393320 556860 393372 556912
rect 425980 556860 426032 556912
rect 495440 556860 495492 556912
rect 3516 556792 3568 556844
rect 360936 556792 360988 556844
rect 370918 556792 370970 556844
rect 462504 556792 462556 556844
rect 207020 556724 207072 556776
rect 248558 556724 248610 556776
rect 333566 556724 333618 556776
rect 461124 556724 461176 556776
rect 218060 556656 218112 556708
rect 321652 556656 321704 556708
rect 332508 556656 332560 556708
rect 462596 556656 462648 556708
rect 227628 556588 227680 556640
rect 269488 556588 269540 556640
rect 312636 556588 312688 556640
rect 459560 556588 459612 556640
rect 233792 556520 233844 556572
rect 234896 556520 234948 556572
rect 339500 556520 339552 556572
rect 453672 556520 453724 556572
rect 193312 556452 193364 556504
rect 359004 556452 359056 556504
rect 360936 556452 360988 556504
rect 518900 556452 518952 556504
rect 227720 556384 227772 556436
rect 283012 556384 283064 556436
rect 291200 556384 291252 556436
rect 461032 556384 461084 556436
rect 193220 556316 193272 556368
rect 276020 556316 276072 556368
rect 296444 556316 296496 556368
rect 512000 556316 512052 556368
rect 226984 556248 227036 556300
rect 247040 556248 247092 556300
rect 395712 556248 395764 556300
rect 513380 556248 513432 556300
rect 226064 556180 226116 556232
rect 254676 556180 254728 556232
rect 399576 556180 399628 556232
rect 571984 556180 572036 556232
rect 117320 555704 117372 555756
rect 235816 556044 235868 556096
rect 235908 556044 235960 556096
rect 234712 555976 234764 556028
rect 114560 555636 114612 555688
rect 234804 555636 234856 555688
rect 107660 555568 107712 555620
rect 234712 555568 234764 555620
rect 86960 555500 87012 555552
rect 234896 555500 234948 555552
rect 3608 555432 3660 555484
rect 261668 556044 261720 556096
rect 364800 556044 364852 556096
rect 223304 554752 223356 554804
rect 232044 554752 232096 554804
rect 451648 555432 451700 555484
rect 580356 555432 580408 555484
rect 454040 554752 454092 554804
rect 211804 554072 211856 554124
rect 233056 554072 233108 554124
rect 118700 554004 118752 554056
rect 233792 554004 233844 554056
rect 451740 554004 451792 554056
rect 580264 554004 580316 554056
rect 3332 553392 3384 553444
rect 10324 553392 10376 553444
rect 223396 553392 223448 553444
rect 232044 553392 232096 553444
rect 453948 553392 454000 553444
rect 468576 553392 468628 553444
rect 60004 552032 60056 552084
rect 232044 552032 232096 552084
rect 452936 551284 452988 551336
rect 574100 551284 574152 551336
rect 160100 550604 160152 550656
rect 232044 550604 232096 550656
rect 2780 549856 2832 549908
rect 232780 549856 232832 549908
rect 453396 549448 453448 549500
rect 455696 549448 455748 549500
rect 104900 548496 104952 548548
rect 232412 548496 232464 548548
rect 26240 547136 26292 547188
rect 232780 547136 232832 547188
rect 453948 546524 454000 546576
rect 457628 546524 457680 546576
rect 176660 545096 176712 545148
rect 232044 545096 232096 545148
rect 453948 545096 454000 545148
rect 536840 545096 536892 545148
rect 60740 544348 60792 544400
rect 232596 544348 232648 544400
rect 453580 544008 453632 544060
rect 455604 544008 455656 544060
rect 67640 542988 67692 543040
rect 228456 542988 228508 543040
rect 453948 542376 454000 542428
rect 468484 542376 468536 542428
rect 233056 541220 233108 541272
rect 233976 541220 234028 541272
rect 11152 540948 11204 541000
rect 232044 540948 232096 541000
rect 453764 540948 453816 541000
rect 462688 540948 462740 541000
rect 42800 540200 42852 540252
rect 225696 540200 225748 540252
rect 223120 539588 223172 539640
rect 232044 539588 232096 539640
rect 189724 538228 189776 538280
rect 232044 538228 232096 538280
rect 224592 536800 224644 536852
rect 232044 536800 232096 536852
rect 453764 536800 453816 536852
rect 463148 536800 463200 536852
rect 479524 536800 479576 536852
rect 580172 536800 580224 536852
rect 453948 535440 454000 535492
rect 520924 535440 520976 535492
rect 80060 534080 80112 534132
rect 232044 534080 232096 534132
rect 229744 532720 229796 532772
rect 232320 532720 232372 532772
rect 453948 532720 454000 532772
rect 461216 532720 461268 532772
rect 1400 529932 1452 529984
rect 232044 529932 232096 529984
rect 96620 528572 96672 528624
rect 232044 528572 232096 528624
rect 3332 527144 3384 527196
rect 19984 527144 20036 527196
rect 453948 527144 454000 527196
rect 471980 527144 472032 527196
rect 224684 525784 224736 525836
rect 232044 525784 232096 525836
rect 453672 524696 453724 524748
rect 455788 524696 455840 524748
rect 128360 524424 128412 524476
rect 232044 524424 232096 524476
rect 452936 523676 452988 523728
rect 453580 523676 453632 523728
rect 4160 521636 4212 521688
rect 232044 521636 232096 521688
rect 453948 521636 454000 521688
rect 461584 521636 461636 521688
rect 453948 520888 454000 520940
rect 457168 520888 457220 520940
rect 204260 520276 204312 520328
rect 232044 520276 232096 520328
rect 223212 518916 223264 518968
rect 232044 518916 232096 518968
rect 453948 518916 454000 518968
rect 475476 518916 475528 518968
rect 88340 516128 88392 516180
rect 232044 516128 232096 516180
rect 3332 514768 3384 514820
rect 224132 514768 224184 514820
rect 453948 514768 454000 514820
rect 500224 514768 500276 514820
rect 453120 514020 453172 514072
rect 453580 514020 453632 514072
rect 453764 513272 453816 513324
rect 465724 513272 465776 513324
rect 227168 510620 227220 510672
rect 232044 510620 232096 510672
rect 541624 510620 541676 510672
rect 580172 510620 580224 510672
rect 453764 509260 453816 509312
rect 462780 509260 462832 509312
rect 228732 506472 228784 506524
rect 232044 506472 232096 506524
rect 222108 505112 222160 505164
rect 232044 505112 232096 505164
rect 232964 504432 233016 504484
rect 232964 504228 233016 504280
rect 453948 503684 454000 503736
rect 464252 503684 464304 503736
rect 51080 502324 51132 502376
rect 232044 502324 232096 502376
rect 3240 502256 3292 502308
rect 234068 502256 234120 502308
rect 220728 500964 220780 501016
rect 232044 500964 232096 501016
rect 453948 499536 454000 499588
rect 548524 499536 548576 499588
rect 453948 498448 454000 498500
rect 457260 498448 457312 498500
rect 179420 495456 179472 495508
rect 232044 495456 232096 495508
rect 453948 492600 454000 492652
rect 498844 492600 498896 492652
rect 224776 488520 224828 488572
rect 232044 488520 232096 488572
rect 453764 488520 453816 488572
rect 464344 488520 464396 488572
rect 453948 487432 454000 487484
rect 458456 487432 458508 487484
rect 230020 485800 230072 485852
rect 231860 485800 231912 485852
rect 453764 485800 453816 485852
rect 480904 485800 480956 485852
rect 453948 484440 454000 484492
rect 458548 484440 458600 484492
rect 213828 484372 213880 484424
rect 232044 484372 232096 484424
rect 471336 484372 471388 484424
rect 580172 484372 580224 484424
rect 453212 482740 453264 482792
rect 459836 482740 459888 482792
rect 222016 481652 222068 481704
rect 232044 481652 232096 481704
rect 125600 480224 125652 480276
rect 232044 480224 232096 480276
rect 453764 480224 453816 480276
rect 543004 480224 543056 480276
rect 52460 477504 52512 477556
rect 232044 477504 232096 477556
rect 453764 477504 453816 477556
rect 465724 477504 465776 477556
rect 453856 476076 453908 476128
rect 549904 476076 549956 476128
rect 3332 475668 3384 475720
rect 8944 475668 8996 475720
rect 120080 474716 120132 474768
rect 232044 474716 232096 474768
rect 453948 474716 454000 474768
rect 556804 474716 556856 474768
rect 230388 473356 230440 473408
rect 231860 473356 231912 473408
rect 453948 472336 454000 472388
rect 458640 472336 458692 472388
rect 55220 471996 55272 472048
rect 232044 471996 232096 472048
rect 453764 471248 453816 471300
rect 458272 471248 458324 471300
rect 202880 470568 202932 470620
rect 232044 470568 232096 470620
rect 486516 470568 486568 470620
rect 579620 470568 579672 470620
rect 453948 469208 454000 469260
rect 529204 469208 529256 469260
rect 452660 468528 452712 468580
rect 454408 468528 454460 468580
rect 453580 466624 453632 466676
rect 455972 466624 456024 466676
rect 218152 465060 218204 465112
rect 232044 465060 232096 465112
rect 218244 464312 218296 464364
rect 222752 464312 222804 464364
rect 453212 464176 453264 464228
rect 455420 464176 455472 464228
rect 57980 463700 58032 463752
rect 232044 463700 232096 463752
rect 226892 462340 226944 462392
rect 232044 462340 232096 462392
rect 453948 462340 454000 462392
rect 475384 462340 475436 462392
rect 48320 460912 48372 460964
rect 232044 460912 232096 460964
rect 164240 459552 164292 459604
rect 232044 459552 232096 459604
rect 453948 459552 454000 459604
rect 504364 459552 504416 459604
rect 452660 458396 452712 458448
rect 454316 458396 454368 458448
rect 220636 458192 220688 458244
rect 231952 458192 232004 458244
rect 216588 456764 216640 456816
rect 232044 456764 232096 456816
rect 19984 456696 20036 456748
rect 231952 456696 232004 456748
rect 453672 455404 453724 455456
rect 462872 455404 462924 455456
rect 453948 454248 454000 454300
rect 457352 454248 457404 454300
rect 228640 454044 228692 454096
rect 232044 454044 232096 454096
rect 228548 452616 228600 452668
rect 232044 452616 232096 452668
rect 453948 452616 454000 452668
rect 465448 452616 465500 452668
rect 153200 451256 153252 451308
rect 232044 451256 232096 451308
rect 453580 450168 453632 450220
rect 455880 450168 455932 450220
rect 3332 449828 3384 449880
rect 227352 449828 227404 449880
rect 453028 447448 453080 447500
rect 454500 447448 454552 447500
rect 453948 444728 454000 444780
rect 460020 444728 460072 444780
rect 229652 444388 229704 444440
rect 232320 444388 232372 444440
rect 220544 442960 220596 443012
rect 232044 442960 232096 443012
rect 225880 441600 225932 441652
rect 232044 441600 232096 441652
rect 228272 440240 228324 440292
rect 232044 440240 232096 440292
rect 453948 440240 454000 440292
rect 544384 440240 544436 440292
rect 453856 440172 453908 440224
rect 502984 440172 503036 440224
rect 453948 437452 454000 437504
rect 489184 437452 489236 437504
rect 453948 436092 454000 436144
rect 461308 436092 461360 436144
rect 453672 435072 453724 435124
rect 456064 435072 456116 435124
rect 158720 433304 158772 433356
rect 231952 433304 232004 433356
rect 79324 433236 79376 433288
rect 232044 433236 232096 433288
rect 453948 430584 454000 430636
rect 526444 430584 526496 430636
rect 462964 429836 463016 429888
rect 580172 429836 580224 429888
rect 229560 429156 229612 429208
rect 231860 429156 231912 429208
rect 91100 427796 91152 427848
rect 232044 427796 232096 427848
rect 453948 427796 454000 427848
rect 525064 427796 525116 427848
rect 85580 426436 85632 426488
rect 232044 426436 232096 426488
rect 453948 426436 454000 426488
rect 494060 426436 494112 426488
rect 168380 425076 168432 425128
rect 232044 425076 232096 425128
rect 453948 425076 454000 425128
rect 555424 425076 555476 425128
rect 452752 425008 452804 425060
rect 541624 425008 541676 425060
rect 122840 423648 122892 423700
rect 232044 423648 232096 423700
rect 3148 422288 3200 422340
rect 228456 422288 228508 422340
rect 453948 420928 454000 420980
rect 463884 420928 463936 420980
rect 209780 419500 209832 419552
rect 232044 419500 232096 419552
rect 453672 418208 453724 418260
rect 456156 418208 456208 418260
rect 491944 418140 491996 418192
rect 579712 418140 579764 418192
rect 453212 416848 453264 416900
rect 455512 416848 455564 416900
rect 227444 415420 227496 415472
rect 231952 415420 232004 415472
rect 453948 413176 454000 413228
rect 458732 413176 458784 413228
rect 227536 412632 227588 412684
rect 232044 412632 232096 412684
rect 82820 409912 82872 409964
rect 232044 409912 232096 409964
rect 3332 409844 3384 409896
rect 225696 409844 225748 409896
rect 452660 408824 452712 408876
rect 454592 408824 454644 408876
rect 10324 408416 10376 408468
rect 232044 408416 232096 408468
rect 453764 407192 453816 407244
rect 456248 407192 456300 407244
rect 453948 407056 454000 407108
rect 491944 407056 491996 407108
rect 453764 404880 453816 404932
rect 460112 404880 460164 404932
rect 565084 404336 565136 404388
rect 580172 404336 580224 404388
rect 132500 401616 132552 401668
rect 232044 401616 232096 401668
rect 453948 401616 454000 401668
rect 463056 401616 463108 401668
rect 452660 400188 452712 400240
rect 454684 400188 454736 400240
rect 190460 398828 190512 398880
rect 232044 398828 232096 398880
rect 453764 398828 453816 398880
rect 465540 398828 465592 398880
rect 232412 398080 232464 398132
rect 233148 398080 233200 398132
rect 3332 397468 3384 397520
rect 228916 397468 228968 397520
rect 232044 397468 232096 397520
rect 231952 397400 232004 397452
rect 225788 395292 225840 395344
rect 234620 395292 234672 395344
rect 95240 394680 95292 394732
rect 232044 394680 232096 394732
rect 453764 394680 453816 394732
rect 461492 394680 461544 394732
rect 453764 393320 453816 393372
rect 464436 393320 464488 393372
rect 453948 391960 454000 392012
rect 491300 391960 491352 392012
rect 191840 390532 191892 390584
rect 232044 390532 232096 390584
rect 453948 389172 454000 389224
rect 465632 389172 465684 389224
rect 453948 386656 454000 386708
rect 457444 386656 457496 386708
rect 453948 385636 454000 385688
rect 456984 385636 457036 385688
rect 24860 385024 24912 385076
rect 232044 385024 232096 385076
rect 195980 383664 196032 383716
rect 232044 383664 232096 383716
rect 453948 383664 454000 383716
rect 502984 383664 503036 383716
rect 453212 382848 453264 382900
rect 460388 382848 460440 382900
rect 230204 382236 230256 382288
rect 232688 382236 232740 382288
rect 453764 378768 453816 378820
rect 457536 378768 457588 378820
rect 225512 378156 225564 378208
rect 232044 378156 232096 378208
rect 460296 378156 460348 378208
rect 580172 378156 580224 378208
rect 453764 375912 453816 375964
rect 458824 375912 458876 375964
rect 29000 375368 29052 375420
rect 232044 375368 232096 375420
rect 230296 374144 230348 374196
rect 232504 374144 232556 374196
rect 230940 374008 230992 374060
rect 231860 374008 231912 374060
rect 453948 372648 454000 372700
rect 456984 372648 457036 372700
rect 224500 372580 224552 372632
rect 232044 372580 232096 372632
rect 223028 371220 223080 371272
rect 232044 371220 232096 371272
rect 453764 371220 453816 371272
rect 476764 371220 476816 371272
rect 453764 369860 453816 369912
rect 534080 369860 534132 369912
rect 226248 368500 226300 368552
rect 232044 368500 232096 368552
rect 453764 368500 453816 368552
rect 486424 368500 486476 368552
rect 453948 367208 454000 367260
rect 458916 367208 458968 367260
rect 231032 367072 231084 367124
rect 231860 367072 231912 367124
rect 453948 365712 454000 365764
rect 464160 365712 464212 365764
rect 453764 364420 453816 364472
rect 463700 364420 463752 364472
rect 461768 364352 461820 364404
rect 580172 364352 580224 364404
rect 194600 362924 194652 362976
rect 232044 362924 232096 362976
rect 227352 361564 227404 361616
rect 232044 361564 232096 361616
rect 453948 361564 454000 361616
rect 462320 361564 462372 361616
rect 232228 360544 232280 360596
rect 233884 360544 233936 360596
rect 453948 358776 454000 358828
rect 562324 358776 562376 358828
rect 453948 357484 454000 357536
rect 456800 357484 456852 357536
rect 213920 356056 213972 356108
rect 232044 356056 232096 356108
rect 453488 355988 453540 356040
rect 459744 355988 459796 356040
rect 224408 355308 224460 355360
rect 232596 355308 232648 355360
rect 451924 355104 451976 355156
rect 452936 355104 452988 355156
rect 228824 351908 228876 351960
rect 232044 351908 232096 351960
rect 229008 350548 229060 350600
rect 232044 350548 232096 350600
rect 453396 350344 453448 350396
rect 454960 350344 455012 350396
rect 232504 349800 232556 349852
rect 232964 349800 233016 349852
rect 227260 349392 227312 349444
rect 228364 349392 228416 349444
rect 69020 349120 69072 349172
rect 232044 349120 232096 349172
rect 452568 348780 452620 348832
rect 454040 348780 454092 348832
rect 228364 347760 228416 347812
rect 232044 347760 232096 347812
rect 453948 347760 454000 347812
rect 478880 347760 478932 347812
rect 453304 347692 453356 347744
rect 454040 347692 454092 347744
rect 453948 347556 454000 347608
rect 459652 347556 459704 347608
rect 230112 346400 230164 346452
rect 232596 346400 232648 346452
rect 3332 346332 3384 346384
rect 60004 346332 60056 346384
rect 222936 345040 222988 345092
rect 232044 345040 232096 345092
rect 201500 344972 201552 345024
rect 231952 344972 232004 345024
rect 71780 344292 71832 344344
rect 222752 344292 222804 344344
rect 452936 343884 452988 343936
rect 454868 343884 454920 343936
rect 452384 342320 452436 342372
rect 454960 342320 455012 342372
rect 102140 342252 102192 342304
rect 232044 342252 232096 342304
rect 453948 342252 454000 342304
rect 471244 342252 471296 342304
rect 453948 342048 454000 342100
rect 458180 342048 458232 342100
rect 74540 340892 74592 340944
rect 231952 340892 232004 340944
rect 21364 340824 21416 340876
rect 232044 340824 232096 340876
rect 234068 338172 234120 338224
rect 236000 338172 236052 338224
rect 447140 338172 447192 338224
rect 465632 338172 465684 338224
rect 34520 338104 34572 338156
rect 232044 338104 232096 338156
rect 226248 338036 226300 338088
rect 580448 338036 580500 338088
rect 229008 337968 229060 338020
rect 580540 337968 580592 338020
rect 409880 337900 409932 337952
rect 452200 337900 452252 337952
rect 419540 337832 419592 337884
rect 464068 337832 464120 337884
rect 405740 337764 405792 337816
rect 462780 337764 462832 337816
rect 394700 337696 394752 337748
rect 456800 337696 456852 337748
rect 231584 337628 231636 337680
rect 244280 337628 244332 337680
rect 387800 337628 387852 337680
rect 458732 337628 458784 337680
rect 225972 337560 226024 337612
rect 253940 337560 253992 337612
rect 376760 337560 376812 337612
rect 454132 337560 454184 337612
rect 233148 337492 233200 337544
rect 262220 337492 262272 337544
rect 333980 337492 334032 337544
rect 452016 337492 452068 337544
rect 233608 337424 233660 337476
rect 278780 337424 278832 337476
rect 448520 337424 448572 337476
rect 580632 337424 580684 337476
rect 224316 337356 224368 337408
rect 243084 337356 243136 337408
rect 249800 337356 249852 337408
rect 454684 337356 454736 337408
rect 428004 337288 428056 337340
rect 465356 337288 465408 337340
rect 430580 337220 430632 337272
rect 462872 337220 462924 337272
rect 434720 337152 434772 337204
rect 455696 337152 455748 337204
rect 451280 337084 451332 337136
rect 464252 337084 464304 337136
rect 227076 336812 227128 336864
rect 245016 336812 245068 336864
rect 3516 336744 3568 336796
rect 262404 336744 262456 336796
rect 225788 336676 225840 336728
rect 378324 336676 378376 336728
rect 378784 336676 378836 336728
rect 380900 336676 380952 336728
rect 400864 336676 400916 336728
rect 402152 336676 402204 336728
rect 422944 336676 422996 336728
rect 423680 336676 423732 336728
rect 427084 336676 427136 336728
rect 427912 336676 427964 336728
rect 446588 336676 446640 336728
rect 449164 336676 449216 336728
rect 450452 336676 450504 336728
rect 485044 336676 485096 336728
rect 222568 336608 222620 336660
rect 266360 336608 266412 336660
rect 342904 336608 342956 336660
rect 461768 336608 461820 336660
rect 222752 336540 222804 336592
rect 241152 336540 241204 336592
rect 244924 336540 244976 336592
rect 246304 336540 246356 336592
rect 275376 336540 275428 336592
rect 283656 336540 283708 336592
rect 367100 336540 367152 336592
rect 464436 336540 464488 336592
rect 232412 336472 232464 336524
rect 291200 336472 291252 336524
rect 357440 336472 357492 336524
rect 461400 336472 461452 336524
rect 229836 336404 229888 336456
rect 296720 336404 296772 336456
rect 441344 336404 441396 336456
rect 462964 336404 463016 336456
rect 224960 336336 225012 336388
rect 460020 336336 460072 336388
rect 21364 336268 21416 336320
rect 269120 336268 269172 336320
rect 277400 336268 277452 336320
rect 454592 336268 454644 336320
rect 165620 336200 165672 336252
rect 463056 336200 463108 336252
rect 24124 336132 24176 336184
rect 323584 336132 323636 336184
rect 342260 336132 342312 336184
rect 459928 336132 459980 336184
rect 28264 336064 28316 336116
rect 413100 336064 413152 336116
rect 424968 336064 425020 336116
rect 486516 336064 486568 336116
rect 26884 335996 26936 336048
rect 416964 335996 417016 336048
rect 420184 335996 420236 336048
rect 436744 335996 436796 336048
rect 440240 335996 440292 336048
rect 457260 335996 457312 336048
rect 222844 335928 222896 335980
rect 233240 335928 233292 335980
rect 280804 335928 280856 335980
rect 282368 335928 282420 335980
rect 381544 335928 381596 335980
rect 389272 335928 389324 335980
rect 405372 335928 405424 335980
rect 448520 335928 448572 335980
rect 225696 335860 225748 335912
rect 234896 335860 234948 335912
rect 407120 335860 407172 335912
rect 433340 335860 433392 335912
rect 405004 335792 405056 335844
rect 425980 335792 426032 335844
rect 320180 335656 320232 335708
rect 451832 335656 451884 335708
rect 360936 335588 360988 335640
rect 366088 335588 366140 335640
rect 380992 335588 381044 335640
rect 456892 335588 456944 335640
rect 232872 334908 232924 334960
rect 282920 334908 282972 334960
rect 364340 334908 364392 334960
rect 455972 334908 456024 334960
rect 233976 334840 234028 334892
rect 298100 334840 298152 334892
rect 340880 334840 340932 334892
rect 452108 334840 452160 334892
rect 230940 334772 230992 334824
rect 375380 334772 375432 334824
rect 415400 334772 415452 334824
rect 451740 334772 451792 334824
rect 234620 334704 234672 334756
rect 241520 334704 241572 334756
rect 259644 334704 259696 334756
rect 452660 334704 452712 334756
rect 232136 334636 232188 334688
rect 438860 334636 438912 334688
rect 44180 334568 44232 334620
rect 453488 334568 453540 334620
rect 23480 333888 23532 333940
rect 324872 333888 324924 333940
rect 398748 333888 398800 333940
rect 565084 333888 565136 333940
rect 286876 333820 286928 333872
rect 471336 333820 471388 333872
rect 131764 333752 131816 333804
rect 397276 333752 397328 333804
rect 418160 333752 418212 333804
rect 462688 333752 462740 333804
rect 255228 333684 255280 333736
rect 477500 333684 477552 333736
rect 253388 333616 253440 333668
rect 460296 333616 460348 333668
rect 275284 333548 275336 333600
rect 479524 333548 479576 333600
rect 157984 333480 158036 333532
rect 356060 333480 356112 333532
rect 374000 333480 374052 333532
rect 451648 333480 451700 333532
rect 225512 333412 225564 333464
rect 231860 333412 231912 333464
rect 248420 333412 248472 333464
rect 465264 333412 465316 333464
rect 201500 333344 201552 333396
rect 457444 333344 457496 333396
rect 200120 333276 200172 333328
rect 462320 333276 462372 333328
rect 129740 333208 129792 333260
rect 458180 333208 458232 333260
rect 224132 333140 224184 333192
rect 390560 333140 390612 333192
rect 429200 333140 429252 333192
rect 463700 333140 463752 333192
rect 40040 333072 40092 333124
rect 311992 333072 312044 333124
rect 347780 333072 347832 333124
rect 452292 333072 452344 333124
rect 352012 333004 352064 333056
rect 451556 333004 451608 333056
rect 234804 331984 234856 332036
rect 271880 331984 271932 332036
rect 232780 331916 232832 331968
rect 303620 331916 303672 331968
rect 307760 331916 307812 331968
rect 456248 331916 456300 331968
rect 267832 331848 267884 331900
rect 453028 331848 453080 331900
rect 231308 330624 231360 330676
rect 317512 330624 317564 330676
rect 349160 330624 349212 330676
rect 454500 330624 454552 330676
rect 233700 330556 233752 330608
rect 281540 330556 281592 330608
rect 311900 330556 311952 330608
rect 455788 330556 455840 330608
rect 231676 330488 231728 330540
rect 382280 330488 382332 330540
rect 270592 330420 270644 330472
rect 271420 330420 271472 330472
rect 346400 330420 346452 330472
rect 347412 330420 347464 330472
rect 228916 329060 228968 329112
rect 400220 329060 400272 329112
rect 284300 327768 284352 327820
rect 455604 327768 455656 327820
rect 183560 327700 183612 327752
rect 454408 327700 454460 327752
rect 394792 326748 394844 326800
rect 395712 326748 395764 326800
rect 233884 326476 233936 326528
rect 383660 326476 383712 326528
rect 251180 326408 251232 326460
rect 453764 326408 453816 326460
rect 223580 326340 223632 326392
rect 456156 326340 456208 326392
rect 329840 325592 329892 325644
rect 580172 325592 580224 325644
rect 231400 325116 231452 325168
rect 353300 325116 353352 325168
rect 229652 325048 229704 325100
rect 477500 325048 477552 325100
rect 184940 324980 184992 325032
rect 449900 324980 449952 325032
rect 121460 324912 121512 324964
rect 457352 324912 457404 324964
rect 233792 323620 233844 323672
rect 346492 323620 346544 323672
rect 228548 323552 228600 323604
rect 280160 323552 280212 323604
rect 292580 323552 292632 323604
rect 454224 323552 454276 323604
rect 340972 322260 341024 322312
rect 457168 322260 457220 322312
rect 81440 322192 81492 322244
rect 225696 322192 225748 322244
rect 229744 322192 229796 322244
rect 420920 322192 420972 322244
rect 231124 320832 231176 320884
rect 510620 320832 510672 320884
rect 3516 320084 3568 320136
rect 220176 320084 220228 320136
rect 231032 319540 231084 319592
rect 310520 319540 310572 319592
rect 229560 319472 229612 319524
rect 393412 319472 393464 319524
rect 78680 319404 78732 319456
rect 453212 319404 453264 319456
rect 228640 318044 228692 318096
rect 276020 318044 276072 318096
rect 284392 318044 284444 318096
rect 454316 318044 454368 318096
rect 387248 316684 387300 316736
rect 568580 316684 568632 316736
rect 260840 315324 260892 315376
rect 449164 315324 449216 315376
rect 189080 315256 189132 315308
rect 448520 315256 448572 315308
rect 556804 313216 556856 313268
rect 580172 313216 580224 313268
rect 49700 312536 49752 312588
rect 458640 312536 458692 312588
rect 345020 309816 345072 309868
rect 437480 309816 437532 309868
rect 329840 309748 329892 309800
rect 457628 309748 457680 309800
rect 369860 308456 369912 308508
rect 436100 308456 436152 308508
rect 198740 308388 198792 308440
rect 453120 308388 453172 308440
rect 216680 307028 216732 307080
rect 456064 307028 456116 307080
rect 3516 306280 3568 306332
rect 317604 306280 317656 306332
rect 324320 305668 324372 305720
rect 374092 305668 374144 305720
rect 389180 305668 389232 305720
rect 400312 305668 400364 305720
rect 433432 305668 433484 305720
rect 547880 305668 547932 305720
rect 234160 305600 234212 305652
rect 498200 305600 498252 305652
rect 345112 303016 345164 303068
rect 402980 303016 403032 303068
rect 150440 302948 150492 303000
rect 346584 302948 346636 303000
rect 394884 302948 394936 303000
rect 533344 302948 533396 303000
rect 115940 302880 115992 302932
rect 458548 302880 458600 302932
rect 234344 301452 234396 301504
rect 580632 301452 580684 301504
rect 103520 300160 103572 300212
rect 259552 300160 259604 300212
rect 232688 300092 232740 300144
rect 408592 300092 408644 300144
rect 468576 299412 468628 299464
rect 580172 299412 580224 299464
rect 173900 297372 173952 297424
rect 455880 297372 455932 297424
rect 228732 296012 228784 296064
rect 322940 296012 322992 296064
rect 309140 295944 309192 295996
rect 484400 295944 484452 295996
rect 284484 294652 284536 294704
rect 502340 294652 502392 294704
rect 84200 294584 84252 294636
rect 458456 294584 458508 294636
rect 3516 293904 3568 293956
rect 461216 293904 461268 293956
rect 231492 291864 231544 291916
rect 335452 291864 335504 291916
rect 9680 291796 9732 291848
rect 251272 291796 251324 291848
rect 320272 291796 320324 291848
rect 556252 291796 556304 291848
rect 59360 290504 59412 290556
rect 242992 290504 243044 290556
rect 231216 290436 231268 290488
rect 516140 290436 516192 290488
rect 172520 289076 172572 289128
rect 438952 289076 439004 289128
rect 147680 284928 147732 284980
rect 341064 284928 341116 284980
rect 361580 284928 361632 284980
rect 549260 284928 549312 284980
rect 316132 282140 316184 282192
rect 378140 282140 378192 282192
rect 144920 280780 144972 280832
rect 280252 280780 280304 280832
rect 292672 280780 292724 280832
rect 396080 280780 396132 280832
rect 234528 273164 234580 273216
rect 580172 273164 580224 273216
rect 53840 272484 53892 272536
rect 255320 272484 255372 272536
rect 313280 272484 313332 272536
rect 567844 272484 567896 272536
rect 226340 269764 226392 269816
rect 385132 269764 385184 269816
rect 369952 268404 370004 268456
rect 467840 268404 467892 268456
rect 135352 268336 135404 268388
rect 375472 268336 375524 268388
rect 3516 267656 3568 267708
rect 461492 267656 461544 267708
rect 294052 262964 294104 263016
rect 427084 262964 427136 263016
rect 142160 262828 142212 262880
rect 293960 262828 294012 262880
rect 151820 257320 151872 257372
rect 328460 257320 328512 257372
rect 227168 255960 227220 256012
rect 411260 255960 411312 256012
rect 3148 255212 3200 255264
rect 459836 255212 459888 255264
rect 226892 254532 226944 254584
rect 422392 254532 422444 254584
rect 89720 250452 89772 250504
rect 422944 250452 422996 250504
rect 100760 247664 100812 247716
rect 360200 247664 360252 247716
rect 33140 246304 33192 246356
rect 306380 246304 306432 246356
rect 225880 245556 225932 245608
rect 580172 245556 580224 245608
rect 66260 239368 66312 239420
rect 458272 239368 458324 239420
rect 70400 235220 70452 235272
rect 382464 235220 382516 235272
rect 230020 233928 230072 233980
rect 386420 233928 386472 233980
rect 13820 233860 13872 233912
rect 405832 233860 405884 233912
rect 99380 232500 99432 232552
rect 278872 232500 278924 232552
rect 3332 215228 3384 215280
rect 447232 215228 447284 215280
rect 376852 206932 376904 206984
rect 579988 206932 580040 206984
rect 3424 202784 3476 202836
rect 461308 202784 461360 202836
rect 475476 193128 475528 193180
rect 580172 193128 580224 193180
rect 3424 188980 3476 189032
rect 464160 188980 464212 189032
rect 208400 180072 208452 180124
rect 452844 180072 452896 180124
rect 247040 179324 247092 179376
rect 580172 179324 580224 179376
rect 169760 174496 169812 174548
rect 455512 174496 455564 174548
rect 233056 173136 233108 173188
rect 423680 173136 423732 173188
rect 224592 166948 224644 167000
rect 580172 166948 580224 167000
rect 211160 164840 211212 164892
rect 431960 164840 432012 164892
rect 3240 164160 3292 164212
rect 211804 164160 211856 164212
rect 35992 157972 36044 158024
rect 244924 157972 244976 158024
rect 527824 153144 527876 153196
rect 579988 153144 580040 153196
rect 300860 152464 300912 152516
rect 527180 152464 527232 152516
rect 3424 150356 3476 150408
rect 385040 150356 385092 150408
rect 62120 145528 62172 145580
rect 275284 145528 275336 145580
rect 287060 139340 287112 139392
rect 580172 139340 580224 139392
rect 469864 138660 469916 138712
rect 580264 138660 580316 138712
rect 263600 123428 263652 123480
rect 331312 123428 331364 123480
rect 3424 111732 3476 111784
rect 206284 111732 206336 111784
rect 480904 100648 480956 100700
rect 580172 100648 580224 100700
rect 3424 97928 3476 97980
rect 267924 97928 267976 97980
rect 295340 91740 295392 91792
rect 474740 91740 474792 91792
rect 30380 90312 30432 90364
rect 343640 90312 343692 90364
rect 209872 87592 209924 87644
rect 452752 87592 452804 87644
rect 224684 86912 224736 86964
rect 580172 86912 580224 86964
rect 231768 86232 231820 86284
rect 365720 86232 365772 86284
rect 3148 85484 3200 85536
rect 199384 85484 199436 85536
rect 232320 80656 232372 80708
rect 416780 80656 416832 80708
rect 223120 73108 223172 73160
rect 580172 73108 580224 73160
rect 3424 71680 3476 71732
rect 200764 71680 200816 71732
rect 77300 69640 77352 69692
rect 378784 69640 378836 69692
rect 85672 65492 85724 65544
rect 360844 65492 360896 65544
rect 69112 64132 69164 64184
rect 383752 64132 383804 64184
rect 227444 59984 227496 60036
rect 397460 59984 397512 60036
rect 241612 57196 241664 57248
rect 368572 57196 368624 57248
rect 149060 55836 149112 55888
rect 405004 55836 405056 55888
rect 287060 54476 287112 54528
rect 434812 54476 434864 54528
rect 27620 51756 27672 51808
rect 269304 51756 269356 51808
rect 269212 51688 269264 51740
rect 400864 51688 400916 51740
rect 321560 47608 321612 47660
rect 528560 47608 528612 47660
rect 234620 47540 234672 47592
rect 455420 47540 455472 47592
rect 507124 46860 507176 46912
rect 580172 46860 580224 46912
rect 334072 46180 334124 46232
rect 489920 46180 489972 46232
rect 3424 45500 3476 45552
rect 338120 45500 338172 45552
rect 298192 43392 298244 43444
rect 470600 43392 470652 43444
rect 398932 39312 398984 39364
rect 459652 39312 459704 39364
rect 40040 35164 40092 35216
rect 453672 35164 453724 35216
rect 3516 33056 3568 33108
rect 456984 33056 457036 33108
rect 474004 33056 474056 33108
rect 580172 33056 580224 33108
rect 237472 32376 237524 32428
rect 372712 32376 372764 32428
rect 228272 31016 228324 31068
rect 332692 31016 332744 31068
rect 489184 31016 489236 31068
rect 506480 31016 506532 31068
rect 276112 29588 276164 29640
rect 488540 29588 488592 29640
rect 143632 28228 143684 28280
rect 353392 28228 353444 28280
rect 226432 25576 226484 25628
rect 336740 25576 336792 25628
rect 230204 25508 230256 25560
rect 343640 25508 343692 25560
rect 368480 25508 368532 25560
rect 538220 25508 538272 25560
rect 161480 24080 161532 24132
rect 379612 24080 379664 24132
rect 394792 24080 394844 24132
rect 514760 24080 514812 24132
rect 3516 22720 3568 22772
rect 189724 22720 189776 22772
rect 325700 22720 325752 22772
rect 473452 22720 473504 22772
rect 168472 21360 168524 21412
rect 307944 21360 307996 21412
rect 3424 20612 3476 20664
rect 288440 20612 288492 20664
rect 538864 20612 538916 20664
rect 579988 20612 580040 20664
rect 421012 18572 421064 18624
rect 463976 18572 464028 18624
rect 367192 17212 367244 17264
rect 392032 17212 392084 17264
rect 418252 17212 418304 17264
rect 444472 17212 444524 17264
rect 371240 15852 371292 15904
rect 533252 15852 533304 15904
rect 307852 14424 307904 14476
rect 326344 14424 326396 14476
rect 465724 14424 465776 14476
rect 509608 14424 509660 14476
rect 230388 13132 230440 13184
rect 273352 13132 273404 13184
rect 110512 13064 110564 13116
rect 167644 13064 167696 13116
rect 235816 13064 235868 13116
rect 314660 13064 314712 13116
rect 357532 13064 357584 13116
rect 544384 13064 544436 13116
rect 126980 11772 127032 11824
rect 128176 11772 128228 11824
rect 184940 11772 184992 11824
rect 186136 11772 186188 11824
rect 109040 11704 109092 11756
rect 217324 11704 217376 11756
rect 227444 11704 227496 11756
rect 227628 11704 227680 11756
rect 270592 11704 270644 11756
rect 526168 11704 526220 11756
rect 77392 10276 77444 10328
rect 220084 10276 220136 10328
rect 221096 10276 221148 10328
rect 327080 10276 327132 10328
rect 331220 10276 331272 10328
rect 515496 10276 515548 10328
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 464344 9596 464396 9648
rect 465172 9596 465224 9648
rect 224868 9188 224920 9240
rect 300768 9188 300820 9240
rect 228824 9120 228876 9172
rect 362316 9120 362368 9172
rect 230296 9052 230348 9104
rect 400128 9052 400180 9104
rect 73804 8984 73856 9036
rect 224224 8984 224276 9036
rect 264980 8984 265032 9036
rect 461676 8984 461728 9036
rect 222936 8916 222988 8968
rect 426164 8916 426216 8968
rect 468484 8916 468536 8968
rect 491116 8916 491168 8968
rect 502984 8916 503036 8968
rect 520740 8916 520792 8968
rect 526444 8916 526496 8968
rect 540796 8916 540848 8968
rect 273260 7964 273312 8016
rect 301964 7964 302016 8016
rect 167184 7896 167236 7948
rect 346400 7896 346452 7948
rect 112812 7828 112864 7880
rect 305000 7828 305052 7880
rect 305552 7828 305604 7880
rect 441712 7828 441764 7880
rect 291292 7760 291344 7812
rect 507676 7760 507728 7812
rect 177856 7692 177908 7744
rect 415492 7692 415544 7744
rect 277492 7624 277544 7676
rect 543188 7624 543240 7676
rect 151912 7556 151964 7608
rect 443000 7556 443052 7608
rect 549904 7556 549956 7608
rect 562048 7556 562100 7608
rect 543004 6876 543056 6928
rect 547880 6876 547932 6928
rect 222016 6808 222068 6860
rect 306748 6808 306800 6860
rect 461584 6808 461636 6860
rect 580172 6808 580224 6860
rect 227352 6740 227404 6792
rect 313832 6740 313884 6792
rect 247592 6672 247644 6724
rect 339500 6672 339552 6724
rect 206192 6604 206244 6656
rect 299480 6604 299532 6656
rect 220728 6536 220780 6588
rect 324412 6536 324464 6588
rect 354680 6536 354732 6588
rect 385960 6536 386012 6588
rect 229836 6468 229888 6520
rect 335360 6468 335412 6520
rect 357532 6468 357584 6520
rect 408500 6468 408552 6520
rect 216588 6400 216640 6452
rect 363512 6400 363564 6452
rect 375288 6400 375340 6452
rect 391940 6400 391992 6452
rect 131764 6332 131816 6384
rect 296812 6332 296864 6384
rect 302332 6332 302384 6384
rect 322112 6332 322164 6384
rect 361120 6332 361172 6384
rect 429292 6332 429344 6384
rect 220544 6264 220596 6316
rect 255872 6264 255924 6316
rect 258264 6264 258316 6316
rect 430672 6264 430724 6316
rect 224500 6196 224552 6248
rect 407212 6196 407264 6248
rect 134156 6128 134208 6180
rect 393320 6128 393372 6180
rect 220636 6060 220688 6112
rect 296076 6060 296128 6112
rect 223488 5992 223540 6044
rect 276020 5992 276072 6044
rect 223028 5924 223080 5976
rect 252376 5924 252428 5976
rect 256700 5924 256752 5976
rect 293684 5924 293736 5976
rect 436744 5516 436796 5568
rect 443828 5516 443880 5568
rect 227444 5380 227496 5432
rect 227628 5380 227680 5432
rect 339868 5176 339920 5228
rect 350540 5176 350592 5228
rect 238852 5108 238904 5160
rect 274824 5108 274876 5160
rect 307944 5108 307996 5160
rect 356060 5108 356112 5160
rect 220452 5040 220504 5092
rect 258080 5040 258132 5092
rect 286600 5040 286652 5092
rect 358912 5040 358964 5092
rect 202696 4972 202748 5024
rect 248512 4972 248564 5024
rect 257068 4972 257120 5024
rect 332600 4972 332652 5024
rect 347872 4972 347924 5024
rect 402520 4972 402572 5024
rect 236092 4904 236144 4956
rect 317328 4904 317380 4956
rect 338672 4904 338724 4956
rect 409972 4904 410024 4956
rect 53748 4836 53800 4888
rect 240232 4836 240284 4888
rect 253480 4836 253532 4888
rect 407304 4836 407356 4888
rect 414020 4836 414072 4888
rect 432052 4836 432104 4888
rect 140044 4768 140096 4820
rect 372620 4768 372672 4820
rect 413100 4768 413152 4820
rect 444380 4768 444432 4820
rect 476764 4768 476816 4820
rect 499396 4768 499448 4820
rect 223396 4020 223448 4072
rect 422300 4156 422352 4208
rect 423772 4156 423824 4208
rect 544476 4156 544528 4208
rect 545488 4156 545540 4208
rect 264152 4088 264204 4140
rect 434444 4088 434496 4140
rect 462412 4088 462464 4140
rect 475384 4088 475436 4140
rect 475936 4088 475988 4140
rect 227536 4020 227588 4072
rect 288992 4020 289044 4072
rect 427268 4020 427320 4072
rect 459560 4020 459612 4072
rect 227260 3952 227312 4004
rect 290188 3952 290240 4004
rect 414296 3952 414348 4004
rect 461032 3952 461084 4004
rect 225420 3884 225472 3936
rect 227352 3884 227404 3936
rect 227720 3884 227772 3936
rect 299664 3884 299716 3936
rect 416688 3884 416740 3936
rect 463884 3884 463936 3936
rect 226156 3816 226208 3868
rect 332600 3816 332652 3868
rect 367836 3816 367888 3868
rect 459192 3816 459244 3868
rect 135260 3748 135312 3800
rect 136456 3748 136508 3800
rect 151820 3748 151872 3800
rect 153016 3748 153068 3800
rect 193220 3748 193272 3800
rect 194416 3748 194468 3800
rect 226340 3748 226392 3800
rect 227536 3748 227588 3800
rect 227628 3748 227680 3800
rect 371700 3748 371752 3800
rect 404820 3748 404872 3800
rect 459744 3748 459796 3800
rect 525064 3748 525116 3800
rect 557356 3748 557408 3800
rect 103336 3680 103388 3732
rect 249892 3680 249944 3732
rect 265348 3680 265400 3732
rect 450544 3680 450596 3732
rect 455696 3680 455748 3732
rect 462596 3680 462648 3732
rect 500224 3680 500276 3732
rect 532516 3680 532568 3732
rect 533344 3680 533396 3732
rect 536104 3680 536156 3732
rect 114008 3612 114060 3664
rect 351920 3612 351972 3664
rect 355232 3612 355284 3664
rect 460940 3612 460992 3664
rect 504364 3612 504416 3664
rect 539600 3612 539652 3664
rect 555424 3612 555476 3664
rect 565636 3612 565688 3664
rect 24216 3544 24268 3596
rect 280804 3544 280856 3596
rect 315028 3544 315080 3596
rect 446404 3544 446456 3596
rect 447784 3544 447836 3596
rect 448612 3544 448664 3596
rect 453304 3544 453356 3596
rect 461124 3544 461176 3596
rect 471244 3544 471296 3596
rect 486424 3544 486476 3596
rect 486516 3544 486568 3596
rect 500592 3544 500644 3596
rect 520924 3544 520976 3596
rect 563244 3544 563296 3596
rect 2780 3476 2832 3528
rect 3700 3476 3752 3528
rect 11060 3476 11112 3528
rect 11980 3476 12032 3528
rect 13544 3476 13596 3528
rect 21364 3476 21416 3528
rect 28908 3476 28960 3528
rect 317420 3476 317472 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 332692 3476 332744 3528
rect 333888 3476 333940 3528
rect 340880 3476 340932 3528
rect 342168 3476 342220 3528
rect 350448 3476 350500 3528
rect 453580 3476 453632 3528
rect 456892 3476 456944 3528
rect 458088 3476 458140 3528
rect 460204 3476 460256 3528
rect 546684 3476 546736 3528
rect 562324 3476 562376 3528
rect 576308 3476 576360 3528
rect 18236 3408 18288 3460
rect 26884 3408 26936 3460
rect 44180 3408 44232 3460
rect 45100 3408 45152 3460
rect 69020 3408 69072 3460
rect 69940 3408 69992 3460
rect 77300 3408 77352 3460
rect 78220 3408 78272 3460
rect 93860 3408 93912 3460
rect 94780 3408 94832 3460
rect 110420 3408 110472 3460
rect 111616 3408 111668 3460
rect 161296 3408 161348 3460
rect 226984 3408 227036 3460
rect 228364 3408 228416 3460
rect 523040 3408 523092 3460
rect 529204 3408 529256 3460
rect 564440 3408 564492 3460
rect 21824 3340 21876 3392
rect 28264 3340 28316 3392
rect 226064 3340 226116 3392
rect 260656 3340 260708 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 365720 3340 365772 3392
rect 367008 3340 367060 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 407120 3340 407172 3392
rect 408408 3340 408460 3392
rect 423680 3340 423732 3392
rect 424968 3340 425020 3392
rect 441528 3340 441580 3392
rect 462504 3340 462556 3392
rect 576124 3340 576176 3392
rect 577412 3340 577464 3392
rect 222108 3272 222160 3324
rect 246396 3272 246448 3324
rect 446404 3272 446456 3324
rect 452384 3272 452436 3324
rect 453580 3272 453632 3324
rect 459008 3272 459060 3324
rect 475936 3272 475988 3324
rect 481732 3272 481784 3324
rect 567844 3272 567896 3324
rect 571524 3272 571576 3324
rect 571984 3272 572036 3324
rect 572720 3272 572772 3324
rect 223212 3204 223264 3256
rect 242900 3204 242952 3256
rect 449808 3204 449860 3256
rect 465080 3204 465132 3256
rect 222752 3136 222804 3188
rect 225604 3136 225656 3188
rect 450912 3136 450964 3188
rect 464528 3136 464580 3188
rect 17040 3068 17092 3120
rect 24124 3068 24176 3120
rect 433248 3068 433300 3120
rect 451924 3068 451976 3120
rect 472624 3000 472676 3052
rect 474556 3000 474608 3052
rect 548524 3000 548576 3052
rect 554964 3000 555016 3052
rect 307760 2864 307812 2916
rect 309048 2864 309100 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 700398 8156 703520
rect 8116 700392 8168 700398
rect 8116 700334 8168 700340
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3422 606112 3478 606121
rect 3422 606047 3478 606056
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3436 577522 3464 606047
rect 21364 579692 21416 579698
rect 21364 579634 21416 579640
rect 3424 577516 3476 577522
rect 3424 577458 3476 577464
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 6920 561808 6972 561814
rect 6920 561750 6972 561756
rect 3424 558204 3476 558210
rect 3424 558146 3476 558152
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2780 549908 2832 549914
rect 2780 549850 2832 549856
rect 1400 529984 1452 529990
rect 1400 529926 1452 529932
rect 18 320784 74 320793
rect 18 320719 74 320728
rect 32 16574 60 320719
rect 32 16546 152 16574
rect 124 354 152 16546
rect 542 354 654 480
rect 124 326 654 354
rect 1412 354 1440 529926
rect 2792 3534 2820 549850
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3344 527202 3372 527847
rect 3332 527196 3384 527202
rect 3332 527138 3384 527144
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3240 502308 3292 502314
rect 3240 502250 3292 502256
rect 3252 501809 3280 502250
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3332 475720 3384 475726
rect 3330 475688 3332 475697
rect 3384 475688 3386 475697
rect 3330 475623 3386 475632
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422346 3188 423535
rect 3148 422340 3200 422346
rect 3148 422282 3200 422288
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3436 241097 3464 558146
rect 3516 556844 3568 556850
rect 3516 556786 3568 556792
rect 3528 371385 3556 556786
rect 3608 555484 3660 555490
rect 3608 555426 3660 555432
rect 3620 462641 3648 555426
rect 4160 521688 4212 521694
rect 4160 521630 4212 521636
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3528 336802 3556 358391
rect 3516 336796 3568 336802
rect 3516 336738 3568 336744
rect 3516 320136 3568 320142
rect 3516 320078 3568 320084
rect 3528 319297 3556 320078
rect 3514 319288 3570 319297
rect 3514 319223 3570 319232
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3516 293956 3568 293962
rect 3516 293898 3568 293904
rect 3528 293185 3556 293898
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 2870 166288 2926 166297
rect 2870 166223 2926 166232
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 166223
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3528 6914 3556 22714
rect 4172 16574 4200 521630
rect 5538 327720 5594 327729
rect 5538 327655 5594 327664
rect 5552 16574 5580 327655
rect 6932 16574 6960 561750
rect 8944 560312 8996 560318
rect 8944 560254 8996 560260
rect 8298 554024 8354 554033
rect 8298 553959 8354 553968
rect 8312 16574 8340 553959
rect 8956 475726 8984 560254
rect 15200 557796 15252 557802
rect 15200 557738 15252 557744
rect 11058 557152 11114 557161
rect 11058 557087 11114 557096
rect 10324 553444 10376 553450
rect 10324 553386 10376 553392
rect 8944 475720 8996 475726
rect 8944 475662 8996 475668
rect 10336 408474 10364 553386
rect 10324 408468 10376 408474
rect 10324 408410 10376 408416
rect 9680 291848 9732 291854
rect 9680 291790 9732 291796
rect 4172 16546 5304 16574
rect 5552 16546 6040 16574
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 3436 6886 3556 6914
rect 3436 6497 3464 6886
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 542 -960 654 326
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 3712 354 3740 3470
rect 5276 480 5304 16546
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 291790
rect 11072 3534 11100 557087
rect 11152 541000 11204 541006
rect 11152 540942 11204 540948
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 540942
rect 13820 233912 13872 233918
rect 13820 233854 13872 233860
rect 13832 16574 13860 233854
rect 15212 16574 15240 557738
rect 19984 527196 20036 527202
rect 19984 527138 20036 527144
rect 19996 456754 20024 527138
rect 19984 456748 20036 456754
rect 19984 456690 20036 456696
rect 21376 340882 21404 579634
rect 21364 340876 21416 340882
rect 21364 340818 21416 340824
rect 21364 336320 21416 336326
rect 21364 336262 21416 336268
rect 19338 333296 19394 333305
rect 19338 333231 19394 333240
rect 19352 16574 19380 333231
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 19352 16546 19472 16574
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11992 354 12020 3470
rect 13556 480 13584 3470
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15948 480 15976 16546
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 17052 480 17080 3062
rect 18248 480 18276 3402
rect 19444 480 19472 16546
rect 21376 3534 21404 336262
rect 23492 333946 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 37278 558240 37334 558249
rect 37278 558175 37334 558184
rect 26240 547188 26292 547194
rect 26240 547130 26292 547136
rect 24860 385076 24912 385082
rect 24860 385018 24912 385024
rect 24124 336184 24176 336190
rect 24124 336126 24176 336132
rect 23480 333940 23532 333946
rect 23480 333882 23532 333888
rect 22098 312488 22154 312497
rect 22098 312423 22154 312432
rect 22112 16574 22140 312423
rect 22112 16546 22600 16574
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21824 3392 21876 3398
rect 20626 3360 20682 3369
rect 21824 3334 21876 3340
rect 20626 3295 20682 3304
rect 20640 480 20668 3295
rect 21836 480 21864 3334
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24136 3126 24164 336126
rect 24872 16574 24900 385018
rect 24872 16546 25360 16574
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 24228 480 24256 3538
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 547130
rect 29000 375420 29052 375426
rect 29000 375362 29052 375368
rect 28264 336116 28316 336122
rect 28264 336058 28316 336064
rect 26884 336048 26936 336054
rect 26884 335990 26936 335996
rect 26896 3466 26924 335990
rect 27620 51808 27672 51814
rect 27620 51750 27672 51756
rect 27632 16574 27660 51750
rect 27632 16546 27752 16574
rect 26884 3460 26936 3466
rect 26884 3402 26936 3408
rect 27724 480 27752 16546
rect 28276 3398 28304 336058
rect 29012 16574 29040 375362
rect 34520 338156 34572 338162
rect 34520 338098 34572 338104
rect 33140 246356 33192 246362
rect 33140 246298 33192 246304
rect 30380 90364 30432 90370
rect 30380 90306 30432 90312
rect 30392 16574 30420 90306
rect 33152 16574 33180 246298
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 33152 16546 33640 16574
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 28920 480 28948 3470
rect 30116 480 30144 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 32402 3496 32458 3505
rect 32402 3431 32458 3440
rect 32416 480 32444 3431
rect 33612 480 33640 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 338098
rect 35898 322144 35954 322153
rect 35898 322079 35954 322088
rect 35912 6914 35940 322079
rect 35992 158024 36044 158030
rect 35992 157966 36044 157972
rect 36004 16574 36032 157966
rect 37292 16574 37320 558175
rect 40052 333130 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 46940 558272 46992 558278
rect 46940 558214 46992 558220
rect 45558 557016 45614 557025
rect 45558 556951 45614 556960
rect 42800 540252 42852 540258
rect 42800 540194 42852 540200
rect 40040 333124 40092 333130
rect 40040 333066 40092 333072
rect 41418 313984 41474 313993
rect 41418 313919 41474 313928
rect 40040 35216 40092 35222
rect 40040 35158 40092 35164
rect 40052 16574 40080 35158
rect 41432 16574 41460 313919
rect 36004 16546 36768 16574
rect 37292 16546 38424 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 35912 6886 36032 6914
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 39578 3632 39634 3641
rect 39578 3567 39634 3576
rect 39592 480 39620 3567
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 540194
rect 44180 334620 44232 334626
rect 44180 334562 44232 334568
rect 44192 3466 44220 334562
rect 44270 316704 44326 316713
rect 44270 316639 44326 316648
rect 44180 3460 44232 3466
rect 44180 3402 44232 3408
rect 44284 480 44312 316639
rect 45572 16574 45600 556951
rect 46952 16574 46980 558214
rect 60004 552084 60056 552090
rect 60004 552026 60056 552032
rect 51080 502376 51132 502382
rect 51080 502318 51132 502324
rect 48320 460964 48372 460970
rect 48320 460906 48372 460912
rect 48332 16574 48360 460906
rect 49700 312588 49752 312594
rect 49700 312530 49752 312536
rect 49712 16574 49740 312530
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 45100 3460 45152 3466
rect 45100 3402 45152 3408
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3402
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 502318
rect 52460 477556 52512 477562
rect 52460 477498 52512 477504
rect 52472 16574 52500 477498
rect 55220 472048 55272 472054
rect 55220 471990 55272 471996
rect 53840 272536 53892 272542
rect 53840 272478 53892 272484
rect 53852 16574 53880 272478
rect 55232 16574 55260 471990
rect 57980 463752 58032 463758
rect 57980 463694 58032 463700
rect 56598 309768 56654 309777
rect 56598 309703 56654 309712
rect 56612 16574 56640 309703
rect 57992 16574 58020 463694
rect 60016 346390 60044 552026
rect 60740 544400 60792 544406
rect 60740 544342 60792 544348
rect 60004 346384 60056 346390
rect 60004 346326 60056 346332
rect 59360 290556 59412 290562
rect 59360 290498 59412 290504
rect 52472 16546 52592 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52564 480 52592 16546
rect 53748 4888 53800 4894
rect 53748 4830 53800 4836
rect 53760 480 53788 4830
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 290498
rect 60752 6914 60780 544342
rect 67640 543040 67692 543046
rect 67640 542982 67692 542988
rect 63498 333432 63554 333441
rect 63498 333367 63554 333376
rect 60830 314120 60886 314129
rect 60830 314055 60886 314064
rect 60844 16574 60872 314055
rect 62120 145580 62172 145586
rect 62120 145522 62172 145528
rect 62132 16574 62160 145522
rect 63512 16574 63540 333367
rect 64878 251832 64934 251841
rect 64878 251767 64934 251776
rect 64892 16574 64920 251767
rect 66260 239420 66312 239426
rect 66260 239362 66312 239368
rect 66272 16574 66300 239362
rect 60844 16546 61608 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 60752 6886 60872 6914
rect 60844 480 60872 6886
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 542982
rect 69020 349172 69072 349178
rect 69020 349114 69072 349120
rect 69032 3466 69060 349114
rect 71792 344350 71820 702986
rect 89180 700330 89208 703520
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 79324 656940 79376 656946
rect 79324 656882 79376 656888
rect 79336 433294 79364 656882
rect 104912 562358 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218256 703582 218836 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 137848 700466 137876 703520
rect 137836 700460 137888 700466
rect 137836 700402 137888 700408
rect 154132 700398 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 157984 700460 158036 700466
rect 157984 700402 158036 700408
rect 131764 700392 131816 700398
rect 131764 700334 131816 700340
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 104900 562352 104952 562358
rect 104900 562294 104952 562300
rect 106280 562216 106332 562222
rect 106280 562158 106332 562164
rect 92480 557864 92532 557870
rect 92480 557806 92532 557812
rect 86960 555552 87012 555558
rect 86960 555494 87012 555500
rect 80060 534132 80112 534138
rect 80060 534074 80112 534080
rect 79324 433288 79376 433294
rect 79324 433230 79376 433236
rect 71780 344344 71832 344350
rect 71780 344286 71832 344292
rect 74540 340944 74592 340950
rect 74540 340886 74592 340892
rect 71778 315344 71834 315353
rect 71778 315279 71834 315288
rect 70400 235272 70452 235278
rect 70400 235214 70452 235220
rect 69112 64184 69164 64190
rect 69112 64126 69164 64132
rect 69020 3460 69072 3466
rect 69020 3402 69072 3408
rect 69124 480 69152 64126
rect 70412 16574 70440 235214
rect 71792 16574 71820 315279
rect 74552 16574 74580 340886
rect 75918 320920 75974 320929
rect 75918 320855 75974 320864
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 74552 16546 75040 16574
rect 69940 3460 69992 3466
rect 69940 3402 69992 3408
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3402
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 73804 9036 73856 9042
rect 73804 8978 73856 8984
rect 73816 480 73844 8978
rect 75012 480 75040 16546
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 320855
rect 78680 319456 78732 319462
rect 78680 319398 78732 319404
rect 77300 69692 77352 69698
rect 77300 69634 77352 69640
rect 77312 3466 77340 69634
rect 78692 16574 78720 319398
rect 80072 16574 80100 534074
rect 85580 426488 85632 426494
rect 85580 426430 85632 426436
rect 82820 409964 82872 409970
rect 82820 409906 82872 409912
rect 81440 322244 81492 322250
rect 81440 322186 81492 322192
rect 81452 16574 81480 322186
rect 82832 16574 82860 409906
rect 84200 294636 84252 294642
rect 84200 294578 84252 294584
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77392 10328 77444 10334
rect 77392 10270 77444 10276
rect 77300 3460 77352 3466
rect 77300 3402 77352 3408
rect 77404 480 77432 10270
rect 78220 3460 78272 3466
rect 78220 3402 78272 3408
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3402
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 294578
rect 85592 6914 85620 426430
rect 85672 65544 85724 65550
rect 85672 65486 85724 65492
rect 85684 16574 85712 65486
rect 86972 16574 87000 555494
rect 88340 516180 88392 516186
rect 88340 516122 88392 516128
rect 88352 16574 88380 516122
rect 91100 427848 91152 427854
rect 91100 427790 91152 427796
rect 89720 250504 89772 250510
rect 89720 250446 89772 250452
rect 89732 16574 89760 250446
rect 91112 16574 91140 427790
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 557806
rect 104900 548548 104952 548554
rect 104900 548490 104952 548496
rect 96620 528624 96672 528630
rect 96620 528566 96672 528572
rect 95240 394732 95292 394738
rect 95240 394674 95292 394680
rect 93858 283520 93914 283529
rect 93858 283455 93914 283464
rect 93872 3466 93900 283455
rect 95252 16574 95280 394674
rect 96632 16574 96660 528566
rect 102140 342304 102192 342310
rect 102140 342246 102192 342252
rect 97998 311128 98054 311137
rect 97998 311063 98054 311072
rect 98012 16574 98040 311063
rect 100760 247716 100812 247722
rect 100760 247658 100812 247664
rect 99380 232552 99432 232558
rect 99380 232494 99432 232500
rect 99392 16574 99420 232494
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93950 15872 94006 15881
rect 93950 15807 94006 15816
rect 93860 3460 93912 3466
rect 93860 3402 93912 3408
rect 93964 480 93992 15807
rect 94780 3460 94832 3466
rect 94780 3402 94832 3408
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3402
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 247658
rect 102152 16574 102180 342246
rect 103520 300212 103572 300218
rect 103520 300154 103572 300160
rect 103532 16574 103560 300154
rect 104912 16574 104940 548490
rect 106292 16574 106320 562158
rect 126980 557592 127032 557598
rect 126980 557534 127032 557540
rect 117320 555756 117372 555762
rect 117320 555698 117372 555704
rect 114560 555688 114612 555694
rect 114560 555630 114612 555636
rect 107660 555620 107712 555626
rect 107660 555562 107712 555568
rect 107672 16574 107700 555562
rect 110418 323640 110474 323649
rect 110418 323575 110474 323584
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102244 480 102272 16546
rect 103336 3732 103388 3738
rect 103336 3674 103388 3680
rect 103348 480 103376 3674
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109040 11756 109092 11762
rect 109040 11698 109092 11704
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 11698
rect 110432 3466 110460 323575
rect 114572 16574 114600 555630
rect 115940 302932 115992 302938
rect 115940 302874 115992 302880
rect 115952 16574 115980 302874
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110512 13116 110564 13122
rect 110512 13058 110564 13064
rect 110420 3460 110472 3466
rect 110420 3402 110472 3408
rect 110524 480 110552 13058
rect 112812 7880 112864 7886
rect 112812 7822 112864 7828
rect 111616 3460 111668 3466
rect 111616 3402 111668 3408
rect 111628 480 111656 3402
rect 112824 480 112852 7822
rect 114008 3664 114060 3670
rect 114008 3606 114060 3612
rect 114020 480 114048 3606
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 555698
rect 118700 554056 118752 554062
rect 118700 553998 118752 554004
rect 118712 6914 118740 553998
rect 125600 480276 125652 480282
rect 125600 480218 125652 480224
rect 120080 474768 120132 474774
rect 120080 474710 120132 474716
rect 118790 296032 118846 296041
rect 118790 295967 118846 295976
rect 118804 16574 118832 295967
rect 120092 16574 120120 474710
rect 122840 423700 122892 423706
rect 122840 423642 122892 423648
rect 121460 324964 121512 324970
rect 121460 324906 121512 324912
rect 121472 16574 121500 324906
rect 122852 16574 122880 423642
rect 124218 333568 124274 333577
rect 124218 333503 124274 333512
rect 124232 16574 124260 333503
rect 118804 16546 119936 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 118712 6886 118832 6914
rect 118804 480 118832 6886
rect 119908 480 119936 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 480218
rect 126992 11830 127020 557534
rect 127072 557048 127124 557054
rect 127072 556990 127124 556996
rect 126980 11824 127032 11830
rect 126980 11766 127032 11772
rect 127084 6914 127112 556990
rect 128360 524476 128412 524482
rect 128360 524418 128412 524424
rect 128372 16574 128400 524418
rect 131776 333810 131804 700334
rect 155960 558340 156012 558346
rect 155960 558282 156012 558288
rect 136640 557932 136692 557938
rect 136640 557874 136692 557880
rect 132500 401668 132552 401674
rect 132500 401610 132552 401616
rect 131764 333804 131816 333810
rect 131764 333746 131816 333752
rect 129740 333260 129792 333266
rect 129740 333202 129792 333208
rect 129752 16574 129780 333202
rect 132512 16574 132540 401610
rect 135258 301472 135314 301481
rect 135258 301407 135314 301416
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 132512 16546 133000 16574
rect 128176 11824 128228 11830
rect 128176 11766 128228 11772
rect 126992 6886 127112 6914
rect 126992 480 127020 6886
rect 128188 480 128216 11766
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 131764 6384 131816 6390
rect 131764 6326 131816 6332
rect 131776 480 131804 6326
rect 132972 480 133000 16546
rect 134156 6180 134208 6186
rect 134156 6122 134208 6128
rect 134168 480 134196 6122
rect 135272 3806 135300 301407
rect 135352 268388 135404 268394
rect 135352 268330 135404 268336
rect 135260 3800 135312 3806
rect 135260 3742 135312 3748
rect 135364 3482 135392 268330
rect 136652 16574 136680 557874
rect 140778 557696 140834 557705
rect 140778 557631 140834 557640
rect 140792 16574 140820 557631
rect 143540 557116 143592 557122
rect 143540 557058 143592 557064
rect 142160 262880 142212 262886
rect 142160 262822 142212 262828
rect 136652 16546 137232 16574
rect 140792 16546 141280 16574
rect 136456 3800 136508 3806
rect 136456 3742 136508 3748
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3742
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 140044 4820 140096 4826
rect 140044 4762 140096 4768
rect 138846 3904 138902 3913
rect 138846 3839 138902 3848
rect 138860 480 138888 3839
rect 140056 480 140084 4762
rect 141252 480 141280 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142172 354 142200 262822
rect 143552 480 143580 557058
rect 153200 451308 153252 451314
rect 153200 451250 153252 451256
rect 146298 336016 146354 336025
rect 146298 335951 146354 335960
rect 144920 280832 144972 280838
rect 144920 280774 144972 280780
rect 143632 28280 143684 28286
rect 143632 28222 143684 28228
rect 143644 16574 143672 28222
rect 144932 16574 144960 280774
rect 146312 16574 146340 335951
rect 150440 303000 150492 303006
rect 150440 302942 150492 302948
rect 147680 284980 147732 284986
rect 147680 284922 147732 284928
rect 147692 16574 147720 284922
rect 149060 55888 149112 55894
rect 149060 55830 149112 55836
rect 149072 16574 149100 55830
rect 150452 16574 150480 302942
rect 151820 257372 151872 257378
rect 151820 257314 151872 257320
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 3806 151860 257314
rect 153212 16574 153240 451250
rect 154578 112432 154634 112441
rect 154578 112367 154634 112376
rect 154592 16574 154620 112367
rect 155972 16574 156000 558282
rect 157338 334656 157394 334665
rect 157338 334591 157394 334600
rect 157352 16574 157380 334591
rect 157996 333538 158024 700402
rect 169772 566506 169800 702406
rect 169760 566500 169812 566506
rect 169760 566442 169812 566448
rect 200764 560924 200816 560930
rect 200764 560866 200816 560872
rect 199384 560584 199436 560590
rect 199384 560526 199436 560532
rect 167644 559360 167696 559366
rect 167644 559302 167696 559308
rect 162860 557660 162912 557666
rect 162860 557602 162912 557608
rect 160100 550656 160152 550662
rect 160100 550598 160152 550604
rect 158720 433356 158772 433362
rect 158720 433298 158772 433304
rect 157984 333532 158036 333538
rect 157984 333474 158036 333480
rect 158732 16574 158760 433298
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 151912 7608 151964 7614
rect 151912 7550 151964 7556
rect 151820 3800 151872 3806
rect 151820 3742 151872 3748
rect 151924 3482 151952 7550
rect 153016 3800 153068 3806
rect 153016 3742 153068 3748
rect 151832 3454 151952 3482
rect 151832 480 151860 3454
rect 153028 480 153056 3742
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 480 160140 550598
rect 161480 24132 161532 24138
rect 161480 24074 161532 24080
rect 161492 16574 161520 24074
rect 162872 16574 162900 557602
rect 164240 459604 164292 459610
rect 164240 459546 164292 459552
rect 164252 16574 164280 459546
rect 165620 336252 165672 336258
rect 165620 336194 165672 336200
rect 165632 16574 165660 336194
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 161296 3460 161348 3466
rect 161296 3402 161348 3408
rect 161308 480 161336 3402
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167656 13122 167684 559302
rect 187700 558000 187752 558006
rect 187700 557942 187752 557948
rect 175280 556912 175332 556918
rect 175280 556854 175332 556860
rect 168380 425128 168432 425134
rect 168380 425070 168432 425076
rect 167644 13116 167696 13122
rect 167644 13058 167696 13064
rect 167184 7948 167236 7954
rect 167184 7890 167236 7896
rect 167196 480 167224 7890
rect 168392 480 168420 425070
rect 171138 336152 171194 336161
rect 171138 336087 171194 336096
rect 169760 174548 169812 174554
rect 169760 174490 169812 174496
rect 168472 21412 168524 21418
rect 168472 21354 168524 21360
rect 168484 16574 168512 21354
rect 169772 16574 169800 174490
rect 171152 16574 171180 336087
rect 173900 297424 173952 297430
rect 173900 297366 173952 297372
rect 172520 289128 172572 289134
rect 172520 289070 172572 289076
rect 172532 16574 172560 289070
rect 168484 16546 169616 16574
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 169588 480 169616 16546
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 297366
rect 175292 16574 175320 556854
rect 176660 545148 176712 545154
rect 176660 545090 176712 545096
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 480 176700 545090
rect 179420 495508 179472 495514
rect 179420 495450 179472 495456
rect 179432 16574 179460 495450
rect 186318 336424 186374 336433
rect 186318 336359 186374 336368
rect 182178 336288 182234 336297
rect 182178 336223 182234 336232
rect 180798 308408 180854 308417
rect 180798 308343 180854 308352
rect 180812 16574 180840 308343
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 177856 7744 177908 7750
rect 177856 7686 177908 7692
rect 177868 480 177896 7686
rect 179050 4040 179106 4049
rect 179050 3975 179106 3984
rect 179064 480 179092 3975
rect 180260 480 180288 16546
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 336223
rect 183560 327752 183612 327758
rect 183560 327694 183612 327700
rect 183572 16574 183600 327694
rect 184940 325032 184992 325038
rect 184940 324974 184992 324980
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11830 184980 324974
rect 186332 16574 186360 336359
rect 187712 16574 187740 557942
rect 197360 557184 197412 557190
rect 197360 557126 197412 557132
rect 193312 556504 193364 556510
rect 193312 556446 193364 556452
rect 193220 556368 193272 556374
rect 193220 556310 193272 556316
rect 189724 538280 189776 538286
rect 189724 538222 189776 538228
rect 189080 315308 189132 315314
rect 189080 315250 189132 315256
rect 189092 16574 189120 315250
rect 189736 22778 189764 538222
rect 190460 398880 190512 398886
rect 190460 398822 190512 398828
rect 189724 22772 189776 22778
rect 189724 22714 189776 22720
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 184940 11824 184992 11830
rect 184940 11766 184992 11772
rect 186136 11824 186188 11830
rect 186136 11766 186188 11772
rect 184938 11656 184994 11665
rect 184938 11591 184994 11600
rect 184952 480 184980 11591
rect 186148 480 186176 11766
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 398822
rect 191840 390584 191892 390590
rect 191840 390526 191892 390532
rect 191852 16574 191880 390526
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 3806 193260 556310
rect 193220 3800 193272 3806
rect 193220 3742 193272 3748
rect 193324 3482 193352 556446
rect 195980 383716 196032 383722
rect 195980 383658 196032 383664
rect 194600 362976 194652 362982
rect 194600 362918 194652 362924
rect 194612 16574 194640 362918
rect 195992 16574 196020 383658
rect 197372 16574 197400 557126
rect 198740 308440 198792 308446
rect 198740 308382 198792 308388
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194416 3800 194468 3806
rect 194416 3742 194468 3748
rect 193232 3454 193352 3482
rect 193232 480 193260 3454
rect 194428 480 194456 3742
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 308382
rect 199396 85542 199424 560526
rect 200120 333328 200172 333334
rect 200120 333270 200172 333276
rect 199384 85536 199436 85542
rect 199384 85478 199436 85484
rect 200132 16574 200160 333270
rect 200776 71738 200804 560866
rect 201512 345030 201540 702986
rect 215300 562488 215352 562494
rect 215300 562430 215352 562436
rect 206284 560720 206336 560726
rect 206284 560662 206336 560668
rect 204260 520328 204312 520334
rect 204260 520270 204312 520276
rect 202880 470620 202932 470626
rect 202880 470562 202932 470568
rect 201500 345024 201552 345030
rect 201500 344966 201552 344972
rect 201500 333396 201552 333402
rect 201500 333338 201552 333344
rect 200764 71732 200816 71738
rect 200764 71674 200816 71680
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 333338
rect 202892 16574 202920 470562
rect 204272 16574 204300 520270
rect 206296 111790 206324 560662
rect 207020 556776 207072 556782
rect 207020 556718 207072 556724
rect 206284 111784 206336 111790
rect 206284 111726 206336 111732
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 202696 5024 202748 5030
rect 202696 4966 202748 4972
rect 202708 480 202736 4966
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206192 6656 206244 6662
rect 206192 6598 206244 6604
rect 206204 480 206232 6598
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 556718
rect 211804 554124 211856 554130
rect 211804 554066 211856 554072
rect 209780 419552 209832 419558
rect 209780 419494 209832 419500
rect 208400 180124 208452 180130
rect 208400 180066 208452 180072
rect 208412 16574 208440 180066
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 9674 209820 419494
rect 211160 164892 211212 164898
rect 211160 164834 211212 164840
rect 209872 87644 209924 87650
rect 209872 87586 209924 87592
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 87586
rect 211172 16574 211200 164834
rect 211816 164218 211844 554066
rect 213828 484424 213880 484430
rect 213828 484366 213880 484372
rect 212538 323776 212594 323785
rect 212538 323711 212594 323720
rect 211804 164212 211856 164218
rect 211804 164154 211856 164160
rect 212552 16574 212580 323711
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 213840 6497 213868 484366
rect 213920 356108 213972 356114
rect 213920 356050 213972 356056
rect 213932 16574 213960 356050
rect 213932 16546 214512 16574
rect 213826 6488 213882 6497
rect 213826 6423 213882 6432
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 562430
rect 217324 559496 217376 559502
rect 217324 559438 217376 559444
rect 216588 456816 216640 456822
rect 216588 456758 216640 456764
rect 216600 6458 216628 456758
rect 216680 307080 216732 307086
rect 216680 307022 216732 307028
rect 216692 16574 216720 307022
rect 216692 16546 216904 16574
rect 216588 6452 216640 6458
rect 216588 6394 216640 6400
rect 216876 480 216904 16546
rect 217336 11762 217364 559438
rect 218060 556708 218112 556714
rect 218060 556650 218112 556656
rect 217324 11756 217376 11762
rect 217324 11698 217376 11704
rect 218072 480 218100 556650
rect 218152 465112 218204 465118
rect 218152 465054 218204 465060
rect 218164 16574 218192 465054
rect 218256 464370 218284 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 227076 700324 227128 700330
rect 227076 700266 227128 700272
rect 233976 700324 234028 700330
rect 233976 700266 234028 700272
rect 224316 562556 224368 562562
rect 224316 562498 224368 562504
rect 220452 562284 220504 562290
rect 220452 562226 220504 562232
rect 220176 560652 220228 560658
rect 220176 560594 220228 560600
rect 220082 559056 220138 559065
rect 220082 558991 220138 559000
rect 218244 464364 218296 464370
rect 218244 464306 218296 464312
rect 218164 16546 219296 16574
rect 219268 480 219296 16546
rect 220096 10334 220124 558991
rect 220188 320142 220216 560594
rect 220464 339017 220492 562226
rect 222844 561060 222896 561066
rect 222844 561002 222896 561008
rect 222108 505164 222160 505170
rect 222108 505106 222160 505112
rect 220728 501016 220780 501022
rect 220728 500958 220780 500964
rect 220636 458244 220688 458250
rect 220636 458186 220688 458192
rect 220544 443012 220596 443018
rect 220544 442954 220596 442960
rect 220450 339008 220506 339017
rect 220450 338943 220506 338952
rect 220176 320136 220228 320142
rect 220176 320078 220228 320084
rect 220084 10328 220136 10334
rect 220084 10270 220136 10276
rect 220556 6322 220584 442954
rect 220544 6316 220596 6322
rect 220544 6258 220596 6264
rect 220648 6118 220676 458186
rect 220740 6594 220768 500958
rect 222016 481704 222068 481710
rect 222016 481646 222068 481652
rect 221096 10328 221148 10334
rect 221096 10270 221148 10276
rect 220728 6588 220780 6594
rect 220728 6530 220780 6536
rect 220636 6112 220688 6118
rect 220636 6054 220688 6060
rect 220452 5092 220504 5098
rect 220452 5034 220504 5040
rect 220464 480 220492 5034
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221108 354 221136 10270
rect 222028 6866 222056 481646
rect 222016 6860 222068 6866
rect 222016 6802 222068 6808
rect 222120 3330 222148 505106
rect 222752 464364 222804 464370
rect 222752 464306 222804 464312
rect 222764 344706 222792 464306
rect 222580 344678 222792 344706
rect 222580 336666 222608 344678
rect 222752 344344 222804 344350
rect 222752 344286 222804 344292
rect 222568 336660 222620 336666
rect 222568 336602 222620 336608
rect 222764 336598 222792 344286
rect 222752 336592 222804 336598
rect 222752 336534 222804 336540
rect 222856 335986 222884 561002
rect 223488 559700 223540 559706
rect 223488 559642 223540 559648
rect 223304 554804 223356 554810
rect 223304 554746 223356 554752
rect 223120 539640 223172 539646
rect 223120 539582 223172 539588
rect 223028 371272 223080 371278
rect 223028 371214 223080 371220
rect 222936 345092 222988 345098
rect 222936 345034 222988 345040
rect 222844 335980 222896 335986
rect 222844 335922 222896 335928
rect 222948 8974 222976 345034
rect 222936 8968 222988 8974
rect 222936 8910 222988 8916
rect 223040 5982 223068 371214
rect 223132 73166 223160 539582
rect 223212 518968 223264 518974
rect 223212 518910 223264 518916
rect 223120 73160 223172 73166
rect 223120 73102 223172 73108
rect 223028 5976 223080 5982
rect 223028 5918 223080 5924
rect 222108 3324 222160 3330
rect 222108 3266 222160 3272
rect 223224 3262 223252 518910
rect 223316 6633 223344 554746
rect 223396 553444 223448 553450
rect 223396 553386 223448 553392
rect 223302 6624 223358 6633
rect 223302 6559 223358 6568
rect 223408 4078 223436 553386
rect 223500 6050 223528 559642
rect 224224 559292 224276 559298
rect 224224 559234 224276 559240
rect 224132 514820 224184 514826
rect 224132 514762 224184 514768
rect 224144 333198 224172 514762
rect 224132 333192 224184 333198
rect 224132 333134 224184 333140
rect 223580 326392 223632 326398
rect 223580 326334 223632 326340
rect 223488 6044 223540 6050
rect 223488 5986 223540 5992
rect 223396 4072 223448 4078
rect 223396 4014 223448 4020
rect 223212 3256 223264 3262
rect 223212 3198 223264 3204
rect 222752 3188 222804 3194
rect 222752 3130 222804 3136
rect 222764 480 222792 3130
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 326334
rect 224236 9042 224264 559234
rect 224328 337414 224356 562498
rect 225972 561876 226024 561882
rect 225972 561818 226024 561824
rect 225694 559600 225750 559609
rect 225694 559535 225750 559544
rect 225604 558476 225656 558482
rect 225604 558418 225656 558424
rect 225420 558408 225472 558414
rect 225420 558350 225472 558356
rect 224866 555928 224922 555937
rect 224866 555863 224922 555872
rect 224592 536852 224644 536858
rect 224592 536794 224644 536800
rect 224500 372632 224552 372638
rect 224500 372574 224552 372580
rect 224408 355360 224460 355366
rect 224408 355302 224460 355308
rect 224316 337408 224368 337414
rect 224316 337350 224368 337356
rect 224224 9036 224276 9042
rect 224224 8978 224276 8984
rect 224420 6225 224448 355302
rect 224512 6254 224540 372574
rect 224604 167006 224632 536794
rect 224684 525836 224736 525842
rect 224684 525778 224736 525784
rect 224592 167000 224644 167006
rect 224592 166942 224644 166948
rect 224696 86970 224724 525778
rect 224776 488572 224828 488578
rect 224776 488514 224828 488520
rect 224684 86964 224736 86970
rect 224684 86906 224736 86912
rect 224500 6248 224552 6254
rect 224406 6216 224462 6225
rect 224500 6190 224552 6196
rect 224406 6151 224462 6160
rect 224788 3777 224816 488514
rect 224880 9246 224908 555863
rect 224960 336388 225012 336394
rect 224960 336330 225012 336336
rect 224972 16574 225000 336330
rect 224972 16546 225184 16574
rect 224868 9240 224920 9246
rect 224868 9182 224920 9188
rect 224774 3768 224830 3777
rect 224774 3703 224830 3712
rect 225156 480 225184 16546
rect 225432 3942 225460 558350
rect 225512 378208 225564 378214
rect 225512 378150 225564 378156
rect 225524 333470 225552 378150
rect 225512 333464 225564 333470
rect 225512 333406 225564 333412
rect 225420 3936 225472 3942
rect 225420 3878 225472 3884
rect 225616 3194 225644 558418
rect 225708 540258 225736 559535
rect 225696 540252 225748 540258
rect 225696 540194 225748 540200
rect 225880 441652 225932 441658
rect 225880 441594 225932 441600
rect 225696 409896 225748 409902
rect 225696 409838 225748 409844
rect 225708 338609 225736 409838
rect 225788 395344 225840 395350
rect 225788 395286 225840 395292
rect 225694 338600 225750 338609
rect 225694 338535 225750 338544
rect 225800 336734 225828 395286
rect 225788 336728 225840 336734
rect 225788 336670 225840 336676
rect 225696 335912 225748 335918
rect 225696 335854 225748 335860
rect 225708 322250 225736 335854
rect 225696 322244 225748 322250
rect 225696 322186 225748 322192
rect 225892 245614 225920 441594
rect 225984 337618 226012 561818
rect 226800 559564 226852 559570
rect 226800 559506 226852 559512
rect 226156 556980 226208 556986
rect 226156 556922 226208 556928
rect 226064 556232 226116 556238
rect 226064 556174 226116 556180
rect 225972 337612 226024 337618
rect 225972 337554 226024 337560
rect 225880 245608 225932 245614
rect 225880 245550 225932 245556
rect 226076 3398 226104 556174
rect 226168 3874 226196 556922
rect 226248 368552 226300 368558
rect 226248 368494 226300 368500
rect 226260 338094 226288 368494
rect 226812 338745 226840 559506
rect 226984 556300 227036 556306
rect 226984 556242 227036 556248
rect 226892 462392 226944 462398
rect 226892 462334 226944 462340
rect 226798 338736 226854 338745
rect 226798 338671 226854 338680
rect 226248 338088 226300 338094
rect 226248 338030 226300 338036
rect 226340 269816 226392 269822
rect 226340 269758 226392 269764
rect 226156 3868 226208 3874
rect 226156 3810 226208 3816
rect 226352 3806 226380 269758
rect 226904 254590 226932 462334
rect 226892 254584 226944 254590
rect 226892 254526 226944 254532
rect 226432 25628 226484 25634
rect 226432 25570 226484 25576
rect 226340 3800 226392 3806
rect 226340 3742 226392 3748
rect 226444 3482 226472 25570
rect 226352 3454 226472 3482
rect 226996 3466 227024 556242
rect 227088 336870 227116 700266
rect 233148 563712 233200 563718
rect 233148 563654 233200 563660
rect 227352 560788 227404 560794
rect 227352 560730 227404 560736
rect 227168 510672 227220 510678
rect 227168 510614 227220 510620
rect 227076 336864 227128 336870
rect 227076 336806 227128 336812
rect 227180 256018 227208 510614
rect 227364 449886 227392 560730
rect 232412 559836 232464 559842
rect 232412 559778 232464 559784
rect 228364 559632 228416 559638
rect 228364 559574 228416 559580
rect 227628 556640 227680 556646
rect 227628 556582 227680 556588
rect 227352 449880 227404 449886
rect 227352 449822 227404 449828
rect 227444 415472 227496 415478
rect 227444 415414 227496 415420
rect 227352 361616 227404 361622
rect 227352 361558 227404 361564
rect 227260 349444 227312 349450
rect 227260 349386 227312 349392
rect 227168 256012 227220 256018
rect 227168 255954 227220 255960
rect 227272 4010 227300 349386
rect 227364 6798 227392 361558
rect 227456 60042 227484 415414
rect 227536 412684 227588 412690
rect 227536 412626 227588 412632
rect 227444 60036 227496 60042
rect 227444 59978 227496 59984
rect 227444 11756 227496 11762
rect 227444 11698 227496 11704
rect 227352 6792 227404 6798
rect 227352 6734 227404 6740
rect 227456 5438 227484 11698
rect 227444 5432 227496 5438
rect 227444 5374 227496 5380
rect 227548 4078 227576 412626
rect 227640 11762 227668 556582
rect 227720 556436 227772 556442
rect 227720 556378 227772 556384
rect 227732 16574 227760 556378
rect 228272 440292 228324 440298
rect 228272 440234 228324 440240
rect 228284 31074 228312 440234
rect 228376 349450 228404 559574
rect 229928 559428 229980 559434
rect 229928 559370 229980 559376
rect 228456 559088 228508 559094
rect 228456 559030 228508 559036
rect 228468 543046 228496 559030
rect 229834 554840 229890 554849
rect 229834 554775 229890 554784
rect 228456 543040 228508 543046
rect 228456 542982 228508 542988
rect 229744 532772 229796 532778
rect 229744 532714 229796 532720
rect 228732 506524 228784 506530
rect 228732 506466 228784 506472
rect 228640 454096 228692 454102
rect 228640 454038 228692 454044
rect 228548 452668 228600 452674
rect 228548 452610 228600 452616
rect 228456 422340 228508 422346
rect 228456 422282 228508 422288
rect 228364 349444 228416 349450
rect 228364 349386 228416 349392
rect 228364 347812 228416 347818
rect 228364 347754 228416 347760
rect 228272 31068 228324 31074
rect 228272 31010 228324 31016
rect 227732 16546 228312 16574
rect 227628 11756 227680 11762
rect 227628 11698 227680 11704
rect 227628 5432 227680 5438
rect 227628 5374 227680 5380
rect 227536 4072 227588 4078
rect 227536 4014 227588 4020
rect 227640 4026 227668 5374
rect 227260 4004 227312 4010
rect 227640 3998 227760 4026
rect 227260 3946 227312 3952
rect 227732 3942 227760 3998
rect 227352 3936 227404 3942
rect 227720 3936 227772 3942
rect 227404 3884 227668 3890
rect 227352 3878 227668 3884
rect 227720 3878 227772 3884
rect 227364 3862 227668 3878
rect 227640 3806 227668 3862
rect 227536 3800 227588 3806
rect 227536 3742 227588 3748
rect 227628 3800 227680 3806
rect 227628 3742 227680 3748
rect 226984 3460 227036 3466
rect 226064 3392 226116 3398
rect 226064 3334 226116 3340
rect 225604 3188 225656 3194
rect 225604 3130 225656 3136
rect 226352 480 226380 3454
rect 226984 3402 227036 3408
rect 227548 480 227576 3742
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228376 3466 228404 347754
rect 228468 339289 228496 422282
rect 228454 339280 228510 339289
rect 228454 339215 228510 339224
rect 228560 323610 228588 452610
rect 228548 323604 228600 323610
rect 228548 323546 228600 323552
rect 228652 318102 228680 454038
rect 228640 318096 228692 318102
rect 228640 318038 228692 318044
rect 228744 296070 228772 506466
rect 229652 444440 229704 444446
rect 229652 444382 229704 444388
rect 229560 429208 229612 429214
rect 229560 429150 229612 429156
rect 228916 397520 228968 397526
rect 228916 397462 228968 397468
rect 228824 351960 228876 351966
rect 228824 351902 228876 351908
rect 228732 296064 228784 296070
rect 228732 296006 228784 296012
rect 228836 9178 228864 351902
rect 228928 329118 228956 397462
rect 229008 350600 229060 350606
rect 229008 350542 229060 350548
rect 229020 338026 229048 350542
rect 229008 338020 229060 338026
rect 229008 337962 229060 337968
rect 228916 329112 228968 329118
rect 228916 329054 228968 329060
rect 229572 319530 229600 429150
rect 229664 325106 229692 444382
rect 229652 325100 229704 325106
rect 229652 325042 229704 325048
rect 229756 322250 229784 532714
rect 229848 336462 229876 554775
rect 229940 338881 229968 559370
rect 232042 555656 232098 555665
rect 232042 555591 232098 555600
rect 232056 554810 232084 555591
rect 232044 554804 232096 554810
rect 232044 554746 232096 554752
rect 232042 554296 232098 554305
rect 232042 554231 232098 554240
rect 232056 553450 232084 554231
rect 232044 553444 232096 553450
rect 232044 553386 232096 553392
rect 232042 552936 232098 552945
rect 232042 552871 232098 552880
rect 232056 552090 232084 552871
rect 232044 552084 232096 552090
rect 232044 552026 232096 552032
rect 232042 551576 232098 551585
rect 232042 551511 232098 551520
rect 232056 550662 232084 551511
rect 232044 550656 232096 550662
rect 232044 550598 232096 550604
rect 231674 548856 231730 548865
rect 231674 548791 231730 548800
rect 231582 509416 231638 509425
rect 231582 509351 231638 509360
rect 230020 485852 230072 485858
rect 230020 485794 230072 485800
rect 229926 338872 229982 338881
rect 229926 338807 229982 338816
rect 229836 336456 229888 336462
rect 229836 336398 229888 336404
rect 229744 322244 229796 322250
rect 229744 322186 229796 322192
rect 229560 319524 229612 319530
rect 229560 319466 229612 319472
rect 230032 233986 230060 485794
rect 231398 479496 231454 479505
rect 231398 479431 231454 479440
rect 231306 476776 231362 476785
rect 231306 476711 231362 476720
rect 230388 473408 230440 473414
rect 230388 473350 230440 473356
rect 230204 382288 230256 382294
rect 230204 382230 230256 382236
rect 230112 346452 230164 346458
rect 230112 346394 230164 346400
rect 230020 233980 230072 233986
rect 230020 233922 230072 233928
rect 228824 9172 228876 9178
rect 228824 9114 228876 9120
rect 229836 6520 229888 6526
rect 229836 6462 229888 6468
rect 228364 3460 228416 3466
rect 228364 3402 228416 3408
rect 229848 480 229876 6462
rect 230124 6361 230152 346394
rect 230216 25566 230244 382230
rect 230296 374196 230348 374202
rect 230296 374138 230348 374144
rect 230204 25560 230256 25566
rect 230204 25502 230256 25508
rect 230308 9110 230336 374138
rect 230400 13190 230428 473350
rect 231214 431896 231270 431905
rect 231214 431831 231270 431840
rect 231122 389736 231178 389745
rect 231122 389671 231178 389680
rect 230940 374060 230992 374066
rect 230940 374002 230992 374008
rect 230952 334830 230980 374002
rect 231032 367124 231084 367130
rect 231032 367066 231084 367072
rect 230940 334824 230992 334830
rect 230940 334766 230992 334772
rect 230478 333160 230534 333169
rect 230478 333095 230534 333104
rect 230492 16574 230520 333095
rect 231044 319598 231072 367066
rect 231136 320890 231164 389671
rect 231124 320884 231176 320890
rect 231124 320826 231176 320832
rect 231032 319592 231084 319598
rect 231032 319534 231084 319540
rect 231228 290494 231256 431831
rect 231320 330682 231348 476711
rect 231308 330676 231360 330682
rect 231308 330618 231360 330624
rect 231412 325174 231440 479431
rect 231490 448896 231546 448905
rect 231490 448831 231546 448840
rect 231400 325168 231452 325174
rect 231400 325110 231452 325116
rect 231504 291922 231532 448831
rect 231596 337686 231624 509351
rect 231584 337680 231636 337686
rect 231584 337622 231636 337628
rect 231688 330546 231716 548791
rect 232424 548554 232452 559778
rect 232686 559736 232742 559745
rect 232686 559671 232742 559680
rect 232594 559464 232650 559473
rect 232594 559399 232650 559408
rect 232502 555248 232558 555257
rect 232502 555183 232558 555192
rect 232412 548548 232464 548554
rect 232412 548490 232464 548496
rect 232042 546136 232098 546145
rect 232042 546071 232098 546080
rect 232056 545154 232084 546071
rect 232044 545148 232096 545154
rect 232044 545090 232096 545096
rect 232042 542056 232098 542065
rect 232042 541991 232098 542000
rect 232056 541006 232084 541991
rect 232044 541000 232096 541006
rect 232044 540942 232096 540948
rect 232042 540016 232098 540025
rect 232042 539951 232098 539960
rect 232056 539646 232084 539951
rect 232044 539640 232096 539646
rect 232044 539582 232096 539588
rect 232042 538656 232098 538665
rect 232042 538591 232098 538600
rect 232056 538286 232084 538591
rect 232044 538280 232096 538286
rect 232044 538222 232096 538228
rect 232042 537296 232098 537305
rect 232042 537231 232098 537240
rect 232056 536858 232084 537231
rect 232044 536852 232096 536858
rect 232044 536794 232096 536800
rect 232042 534576 232098 534585
rect 232042 534511 232098 534520
rect 232056 534138 232084 534511
rect 232044 534132 232096 534138
rect 232044 534074 232096 534080
rect 232318 533216 232374 533225
rect 232318 533151 232374 533160
rect 232332 532778 232360 533151
rect 232320 532772 232372 532778
rect 232320 532714 232372 532720
rect 232042 530496 232098 530505
rect 232042 530431 232098 530440
rect 232056 529990 232084 530431
rect 232044 529984 232096 529990
rect 232044 529926 232096 529932
rect 232042 529136 232098 529145
rect 232042 529071 232098 529080
rect 232056 528630 232084 529071
rect 232044 528624 232096 528630
rect 232044 528566 232096 528572
rect 232042 526416 232098 526425
rect 232042 526351 232098 526360
rect 232056 525842 232084 526351
rect 232044 525836 232096 525842
rect 232044 525778 232096 525784
rect 232042 525056 232098 525065
rect 232042 524991 232098 525000
rect 232056 524482 232084 524991
rect 232044 524476 232096 524482
rect 232044 524418 232096 524424
rect 232042 522336 232098 522345
rect 232042 522271 232098 522280
rect 232056 521694 232084 522271
rect 232044 521688 232096 521694
rect 232044 521630 232096 521636
rect 232044 520328 232096 520334
rect 232042 520296 232044 520305
rect 232096 520296 232098 520305
rect 232042 520231 232098 520240
rect 232044 518968 232096 518974
rect 232042 518936 232044 518945
rect 232096 518936 232098 518945
rect 232042 518871 232098 518880
rect 232042 516216 232098 516225
rect 232042 516151 232044 516160
rect 232096 516151 232098 516160
rect 232044 516122 232096 516128
rect 232042 510776 232098 510785
rect 232042 510711 232098 510720
rect 232056 510678 232084 510711
rect 232044 510672 232096 510678
rect 232044 510614 232096 510620
rect 231766 508056 231822 508065
rect 231766 507991 231822 508000
rect 231676 330540 231728 330546
rect 231676 330482 231728 330488
rect 231492 291916 231544 291922
rect 231492 291858 231544 291864
rect 231216 290488 231268 290494
rect 231216 290430 231268 290436
rect 231780 86290 231808 507991
rect 232042 506696 232098 506705
rect 232042 506631 232098 506640
rect 232056 506530 232084 506631
rect 232044 506524 232096 506530
rect 232044 506466 232096 506472
rect 232042 505336 232098 505345
rect 232042 505271 232098 505280
rect 232056 505170 232084 505271
rect 232044 505164 232096 505170
rect 232044 505106 232096 505112
rect 232042 502616 232098 502625
rect 232042 502551 232098 502560
rect 232056 502382 232084 502551
rect 232044 502376 232096 502382
rect 232044 502318 232096 502324
rect 232042 501256 232098 501265
rect 232042 501191 232098 501200
rect 232056 501022 232084 501191
rect 232044 501016 232096 501022
rect 232044 500958 232096 500964
rect 232042 496496 232098 496505
rect 232042 496431 232098 496440
rect 232056 495514 232084 496431
rect 232044 495508 232096 495514
rect 232044 495450 232096 495456
rect 232042 489696 232098 489705
rect 232042 489631 232098 489640
rect 232056 488578 232084 489631
rect 232044 488572 232096 488578
rect 232044 488514 232096 488520
rect 231858 486976 231914 486985
rect 231858 486911 231914 486920
rect 231872 485858 231900 486911
rect 231860 485852 231912 485858
rect 231860 485794 231912 485800
rect 232042 485616 232098 485625
rect 232042 485551 232098 485560
rect 232056 484430 232084 485551
rect 232044 484424 232096 484430
rect 232044 484366 232096 484372
rect 232042 482896 232098 482905
rect 232042 482831 232098 482840
rect 232056 481710 232084 482831
rect 232044 481704 232096 481710
rect 232044 481646 232096 481652
rect 232042 481536 232098 481545
rect 232042 481471 232098 481480
rect 232056 480282 232084 481471
rect 232044 480276 232096 480282
rect 232044 480218 232096 480224
rect 232042 478136 232098 478145
rect 232042 478071 232098 478080
rect 232056 477562 232084 478071
rect 232044 477556 232096 477562
rect 232044 477498 232096 477504
rect 232042 475416 232098 475425
rect 232042 475351 232098 475360
rect 232056 474774 232084 475351
rect 232044 474768 232096 474774
rect 232044 474710 232096 474716
rect 231858 474056 231914 474065
rect 231858 473991 231914 474000
rect 231872 473414 231900 473991
rect 231860 473408 231912 473414
rect 231860 473350 231912 473356
rect 232042 472696 232098 472705
rect 232042 472631 232098 472640
rect 232056 472054 232084 472631
rect 232044 472048 232096 472054
rect 232044 471990 232096 471996
rect 232042 471336 232098 471345
rect 232042 471271 232098 471280
rect 232056 470626 232084 471271
rect 232044 470620 232096 470626
rect 232044 470562 232096 470568
rect 232042 465896 232098 465905
rect 232042 465831 232098 465840
rect 232056 465118 232084 465831
rect 232044 465112 232096 465118
rect 232044 465054 232096 465060
rect 232042 464536 232098 464545
rect 232042 464471 232098 464480
rect 232056 463758 232084 464471
rect 232044 463752 232096 463758
rect 232044 463694 232096 463700
rect 232042 463176 232098 463185
rect 232042 463111 232098 463120
rect 232056 462398 232084 463111
rect 232044 462392 232096 462398
rect 232044 462334 232096 462340
rect 232042 461816 232098 461825
rect 232042 461751 232098 461760
rect 232056 460970 232084 461751
rect 232044 460964 232096 460970
rect 232044 460906 232096 460912
rect 232042 460456 232098 460465
rect 232042 460391 232098 460400
rect 232056 459610 232084 460391
rect 232044 459604 232096 459610
rect 232044 459546 232096 459552
rect 231950 458416 232006 458425
rect 231950 458351 232006 458360
rect 231964 458250 231992 458351
rect 231952 458244 232004 458250
rect 231952 458186 232004 458192
rect 232042 457056 232098 457065
rect 232042 456991 232098 457000
rect 232056 456822 232084 456991
rect 232044 456816 232096 456822
rect 232044 456758 232096 456764
rect 231952 456748 232004 456754
rect 231952 456690 232004 456696
rect 231964 455705 231992 456690
rect 231950 455696 232006 455705
rect 231950 455631 232006 455640
rect 232042 454336 232098 454345
rect 232042 454271 232098 454280
rect 232056 454102 232084 454271
rect 232044 454096 232096 454102
rect 232044 454038 232096 454044
rect 232042 452976 232098 452985
rect 232042 452911 232098 452920
rect 232056 452674 232084 452911
rect 232044 452668 232096 452674
rect 232044 452610 232096 452616
rect 232042 451616 232098 451625
rect 232042 451551 232098 451560
rect 232056 451314 232084 451551
rect 232044 451308 232096 451314
rect 232044 451250 232096 451256
rect 232318 444816 232374 444825
rect 232318 444751 232374 444760
rect 232332 444446 232360 444751
rect 232320 444440 232372 444446
rect 232320 444382 232372 444388
rect 232042 443456 232098 443465
rect 232042 443391 232098 443400
rect 232056 443018 232084 443391
rect 232044 443012 232096 443018
rect 232044 442954 232096 442960
rect 232042 442096 232098 442105
rect 232042 442031 232098 442040
rect 232056 441658 232084 442031
rect 232044 441652 232096 441658
rect 232044 441594 232096 441600
rect 232042 440736 232098 440745
rect 232042 440671 232098 440680
rect 232056 440298 232084 440671
rect 232044 440292 232096 440298
rect 232044 440234 232096 440240
rect 231950 434616 232006 434625
rect 231950 434551 232006 434560
rect 231964 433362 231992 434551
rect 231952 433356 232004 433362
rect 231952 433298 232004 433304
rect 232044 433288 232096 433294
rect 232042 433256 232044 433265
rect 232096 433256 232098 433265
rect 232042 433191 232098 433200
rect 231858 430536 231914 430545
rect 231858 430471 231914 430480
rect 231872 429214 231900 430471
rect 231860 429208 231912 429214
rect 231860 429150 231912 429156
rect 232042 429176 232098 429185
rect 232042 429111 232098 429120
rect 232056 427854 232084 429111
rect 232044 427848 232096 427854
rect 232044 427790 232096 427796
rect 232044 426488 232096 426494
rect 232042 426456 232044 426465
rect 232096 426456 232098 426465
rect 232042 426391 232098 426400
rect 232044 425128 232096 425134
rect 232042 425096 232044 425105
rect 232096 425096 232098 425105
rect 232042 425031 232098 425040
rect 232042 423736 232098 423745
rect 232042 423671 232044 423680
rect 232096 423671 232098 423680
rect 232044 423642 232096 423648
rect 232042 419656 232098 419665
rect 232042 419591 232098 419600
rect 232056 419558 232084 419591
rect 232044 419552 232096 419558
rect 232044 419494 232096 419500
rect 231950 416256 232006 416265
rect 231950 416191 232006 416200
rect 231964 415478 231992 416191
rect 231952 415472 232004 415478
rect 231952 415414 232004 415420
rect 232042 413536 232098 413545
rect 232042 413471 232098 413480
rect 232056 412690 232084 413471
rect 232044 412684 232096 412690
rect 232044 412626 232096 412632
rect 232042 410816 232098 410825
rect 232042 410751 232098 410760
rect 232056 409970 232084 410751
rect 232044 409964 232096 409970
rect 232044 409906 232096 409912
rect 232044 408468 232096 408474
rect 232044 408410 232096 408416
rect 232056 408105 232084 408410
rect 232042 408096 232098 408105
rect 232042 408031 232098 408040
rect 232410 404016 232466 404025
rect 232410 403951 232466 403960
rect 232042 402656 232098 402665
rect 232042 402591 232098 402600
rect 232056 401674 232084 402591
rect 232044 401668 232096 401674
rect 232044 401610 232096 401616
rect 232042 399936 232098 399945
rect 232042 399871 232098 399880
rect 232056 398886 232084 399871
rect 232044 398880 232096 398886
rect 232044 398822 232096 398828
rect 232424 398138 232452 403951
rect 232412 398132 232464 398138
rect 232412 398074 232464 398080
rect 232042 397896 232098 397905
rect 232042 397831 232098 397840
rect 232056 397526 232084 397831
rect 232044 397520 232096 397526
rect 232044 397462 232096 397468
rect 231952 397452 232004 397458
rect 231952 397394 232004 397400
rect 231964 396545 231992 397394
rect 231950 396536 232006 396545
rect 231950 396471 232006 396480
rect 232042 395176 232098 395185
rect 232042 395111 232098 395120
rect 232056 394738 232084 395111
rect 232044 394732 232096 394738
rect 232044 394674 232096 394680
rect 232410 393816 232466 393825
rect 232410 393751 232466 393760
rect 232042 391096 232098 391105
rect 232042 391031 232098 391040
rect 232056 390590 232084 391031
rect 232044 390584 232096 390590
rect 232044 390526 232096 390532
rect 232042 385656 232098 385665
rect 232042 385591 232098 385600
rect 232056 385082 232084 385591
rect 232044 385076 232096 385082
rect 232044 385018 232096 385024
rect 232042 384296 232098 384305
rect 232042 384231 232098 384240
rect 232056 383722 232084 384231
rect 232044 383716 232096 383722
rect 232044 383658 232096 383664
rect 232042 378856 232098 378865
rect 232042 378791 232098 378800
rect 232056 378214 232084 378791
rect 232044 378208 232096 378214
rect 232044 378150 232096 378156
rect 232134 376816 232190 376825
rect 232134 376751 232190 376760
rect 232042 375456 232098 375465
rect 232042 375391 232044 375400
rect 232096 375391 232098 375400
rect 232044 375362 232096 375368
rect 231858 374096 231914 374105
rect 231858 374031 231860 374040
rect 231912 374031 231914 374040
rect 231860 374002 231912 374008
rect 232042 372736 232098 372745
rect 232042 372671 232098 372680
rect 232056 372638 232084 372671
rect 232044 372632 232096 372638
rect 232044 372574 232096 372580
rect 232042 371376 232098 371385
rect 232042 371311 232098 371320
rect 232056 371278 232084 371311
rect 232044 371272 232096 371278
rect 232044 371214 232096 371220
rect 232042 368656 232098 368665
rect 232042 368591 232098 368600
rect 232056 368558 232084 368591
rect 232044 368552 232096 368558
rect 232044 368494 232096 368500
rect 231858 367296 231914 367305
rect 231858 367231 231914 367240
rect 231872 367130 231900 367231
rect 231860 367124 231912 367130
rect 231860 367066 231912 367072
rect 232042 363216 232098 363225
rect 232042 363151 232098 363160
rect 232056 362982 232084 363151
rect 232044 362976 232096 362982
rect 232044 362918 232096 362924
rect 232042 361856 232098 361865
rect 232042 361791 232098 361800
rect 232056 361622 232084 361791
rect 232044 361616 232096 361622
rect 232044 361558 232096 361564
rect 232042 357096 232098 357105
rect 232042 357031 232098 357040
rect 232056 356114 232084 357031
rect 232044 356108 232096 356114
rect 232044 356050 232096 356056
rect 232042 353016 232098 353025
rect 232042 352951 232098 352960
rect 232056 351966 232084 352951
rect 232044 351960 232096 351966
rect 232044 351902 232096 351908
rect 232042 351656 232098 351665
rect 232042 351591 232098 351600
rect 232056 350606 232084 351591
rect 232044 350600 232096 350606
rect 232044 350542 232096 350548
rect 232042 350296 232098 350305
rect 232042 350231 232098 350240
rect 232056 349178 232084 350231
rect 232044 349172 232096 349178
rect 232044 349114 232096 349120
rect 232042 348936 232098 348945
rect 232042 348871 232098 348880
rect 232056 347818 232084 348871
rect 232044 347812 232096 347818
rect 232044 347754 232096 347760
rect 232042 346216 232098 346225
rect 232042 346151 232098 346160
rect 232056 345098 232084 346151
rect 232044 345092 232096 345098
rect 232044 345034 232096 345040
rect 231952 345024 232004 345030
rect 231952 344966 232004 344972
rect 231964 344865 231992 344966
rect 231950 344856 232006 344865
rect 231950 344791 232006 344800
rect 232042 343496 232098 343505
rect 232042 343431 232098 343440
rect 232056 342310 232084 343431
rect 232044 342304 232096 342310
rect 232044 342246 232096 342252
rect 231950 342136 232006 342145
rect 231950 342071 232006 342080
rect 231964 340950 231992 342071
rect 231952 340944 232004 340950
rect 231952 340886 232004 340892
rect 232044 340876 232096 340882
rect 232044 340818 232096 340824
rect 232056 340785 232084 340818
rect 232042 340776 232098 340785
rect 232042 340711 232098 340720
rect 232042 339416 232098 339425
rect 232042 339351 232098 339360
rect 232056 338162 232084 339351
rect 232044 338156 232096 338162
rect 232044 338098 232096 338104
rect 232148 334694 232176 376751
rect 232228 360596 232280 360602
rect 232228 360538 232280 360544
rect 232240 339969 232268 360538
rect 232318 354376 232374 354385
rect 232318 354311 232374 354320
rect 232226 339960 232282 339969
rect 232226 339895 232282 339904
rect 232136 334688 232188 334694
rect 232136 334630 232188 334636
rect 231860 333464 231912 333470
rect 231860 333406 231912 333412
rect 231768 86284 231820 86290
rect 231768 86226 231820 86232
rect 230492 16546 231072 16574
rect 230388 13184 230440 13190
rect 230388 13126 230440 13132
rect 230296 9104 230348 9110
rect 230296 9046 230348 9052
rect 230110 6352 230166 6361
rect 230110 6287 230166 6296
rect 231044 480 231072 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 228702 -960 228814 326
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 231872 354 231900 333406
rect 232332 80714 232360 354311
rect 232424 336530 232452 393751
rect 232516 374202 232544 555183
rect 232608 544406 232636 559399
rect 232700 547874 232728 559671
rect 232780 558952 232832 558958
rect 232780 558894 232832 558900
rect 232792 549914 232820 558894
rect 232872 558068 232924 558074
rect 232872 558010 232924 558016
rect 232884 557534 232912 558010
rect 232884 557506 233004 557534
rect 232780 549908 232832 549914
rect 232780 549850 232832 549856
rect 232700 547846 232820 547874
rect 232792 547194 232820 547846
rect 232780 547188 232832 547194
rect 232780 547130 232832 547136
rect 232596 544400 232648 544406
rect 232596 544342 232648 544348
rect 232976 504490 233004 557506
rect 233054 556064 233110 556073
rect 233054 555999 233110 556008
rect 233068 554130 233096 555999
rect 233056 554124 233108 554130
rect 233056 554066 233108 554072
rect 233056 541272 233108 541278
rect 233056 541214 233108 541220
rect 232964 504484 233016 504490
rect 232964 504426 233016 504432
rect 233068 504370 233096 541214
rect 232884 504342 233096 504370
rect 232884 493785 232912 504342
rect 232964 504280 233016 504286
rect 232964 504222 233016 504228
rect 232870 493776 232926 493785
rect 232870 493711 232926 493720
rect 232870 450256 232926 450265
rect 232870 450191 232926 450200
rect 232594 435976 232650 435985
rect 232594 435911 232650 435920
rect 232504 374196 232556 374202
rect 232504 374138 232556 374144
rect 232502 364576 232558 364585
rect 232502 364511 232558 364520
rect 232516 354674 232544 364511
rect 232608 355366 232636 435911
rect 232778 422376 232834 422385
rect 232778 422311 232834 422320
rect 232686 382936 232742 382945
rect 232686 382871 232742 382880
rect 232700 382294 232728 382871
rect 232688 382288 232740 382294
rect 232688 382230 232740 382236
rect 232596 355360 232648 355366
rect 232596 355302 232648 355308
rect 232516 354646 232728 354674
rect 232504 349852 232556 349858
rect 232504 349794 232556 349800
rect 232516 339833 232544 349794
rect 232594 347576 232650 347585
rect 232594 347511 232650 347520
rect 232608 346458 232636 347511
rect 232596 346452 232648 346458
rect 232596 346394 232648 346400
rect 232502 339824 232558 339833
rect 232502 339759 232558 339768
rect 232412 336524 232464 336530
rect 232412 336466 232464 336472
rect 232700 300150 232728 354646
rect 232792 331974 232820 422311
rect 232884 334966 232912 450191
rect 232976 349858 233004 504222
rect 233160 495145 233188 563654
rect 233884 558136 233936 558142
rect 233884 558078 233936 558084
rect 233792 556572 233844 556578
rect 233792 556514 233844 556520
rect 233804 554062 233832 556514
rect 233792 554056 233844 554062
rect 233792 553998 233844 554004
rect 233146 495136 233202 495145
rect 233146 495071 233202 495080
rect 233054 412176 233110 412185
rect 233054 412111 233110 412120
rect 232964 349852 233016 349858
rect 232964 349794 233016 349800
rect 232872 334960 232924 334966
rect 232872 334902 232924 334908
rect 232780 331968 232832 331974
rect 232780 331910 232832 331916
rect 232688 300144 232740 300150
rect 232688 300086 232740 300092
rect 233068 173194 233096 412111
rect 233148 398132 233200 398138
rect 233148 398074 233200 398080
rect 233160 337550 233188 398074
rect 233790 380216 233846 380225
rect 233790 380151 233846 380160
rect 233606 359136 233662 359145
rect 233606 359071 233662 359080
rect 233148 337544 233200 337550
rect 233148 337486 233200 337492
rect 233620 337482 233648 359071
rect 233698 355736 233754 355745
rect 233698 355671 233754 355680
rect 233608 337476 233660 337482
rect 233608 337418 233660 337424
rect 233240 335980 233292 335986
rect 233240 335922 233292 335928
rect 233056 173188 233108 173194
rect 233056 173130 233108 173136
rect 232320 80708 232372 80714
rect 232320 80650 232372 80656
rect 233252 16574 233280 335922
rect 233712 330614 233740 355671
rect 233700 330608 233752 330614
rect 233700 330550 233752 330556
rect 233804 323678 233832 380151
rect 233896 360602 233924 558078
rect 233988 541278 234016 700266
rect 234252 572008 234304 572014
rect 234252 571950 234304 571956
rect 234160 570648 234212 570654
rect 234160 570590 234212 570596
rect 234066 555112 234122 555121
rect 234066 555047 234122 555056
rect 233976 541272 234028 541278
rect 233976 541214 234028 541220
rect 234080 502314 234108 555047
rect 234068 502308 234120 502314
rect 234068 502250 234120 502256
rect 234172 484265 234200 570590
rect 234158 484256 234214 484265
rect 234158 484191 234214 484200
rect 234264 468625 234292 571950
rect 234344 563780 234396 563786
rect 234344 563722 234396 563728
rect 234250 468616 234306 468625
rect 234250 468551 234306 468560
rect 234250 438696 234306 438705
rect 234250 438631 234306 438640
rect 234066 421016 234122 421025
rect 234066 420951 234122 420960
rect 233974 392456 234030 392465
rect 233974 392391 234030 392400
rect 233884 360596 233936 360602
rect 233884 360538 233936 360544
rect 233882 360496 233938 360505
rect 233882 360431 233938 360440
rect 233896 326534 233924 360431
rect 233988 334898 234016 392391
rect 234080 338230 234108 420951
rect 234158 401296 234214 401305
rect 234158 401231 234214 401240
rect 234068 338224 234120 338230
rect 234068 338166 234120 338172
rect 233976 334892 234028 334898
rect 233976 334834 234028 334840
rect 233884 326528 233936 326534
rect 233884 326470 233936 326476
rect 233792 323672 233844 323678
rect 233792 323614 233844 323620
rect 234172 305658 234200 401231
rect 234264 338201 234292 438631
rect 234356 409465 234384 563722
rect 234528 562420 234580 562426
rect 234528 562362 234580 562368
rect 234434 555520 234490 555529
rect 234434 555455 234490 555464
rect 234342 409456 234398 409465
rect 234342 409391 234398 409400
rect 234342 405376 234398 405385
rect 234342 405311 234398 405320
rect 234250 338192 234306 338201
rect 234250 338127 234306 338136
rect 234160 305652 234212 305658
rect 234160 305594 234212 305600
rect 234356 301510 234384 405311
rect 234448 358465 234476 555455
rect 234540 547505 234568 562362
rect 234526 547496 234582 547505
rect 234526 547431 234582 547440
rect 234526 499216 234582 499225
rect 234526 499151 234582 499160
rect 234434 358456 234490 358465
rect 234434 358391 234490 358400
rect 234344 301504 234396 301510
rect 234344 301446 234396 301452
rect 234540 273222 234568 499151
rect 234632 395350 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 255320 700460 255372 700466
rect 255320 700402 255372 700408
rect 237380 630692 237432 630698
rect 237380 630634 237432 630640
rect 234896 559904 234948 559910
rect 234896 559846 234948 559852
rect 234712 559768 234764 559774
rect 234712 559710 234764 559716
rect 234724 556322 234752 559710
rect 234802 559192 234858 559201
rect 234802 559127 234858 559136
rect 234816 556458 234844 559127
rect 234908 556578 234936 559846
rect 235816 559156 235868 559162
rect 235816 559098 235868 559104
rect 234896 556572 234948 556578
rect 234896 556514 234948 556520
rect 234816 556430 234936 556458
rect 234724 556294 234844 556322
rect 234712 556028 234764 556034
rect 234712 555970 234764 555976
rect 234724 555626 234752 555970
rect 234816 555694 234844 556294
rect 234804 555688 234856 555694
rect 234804 555630 234856 555636
rect 234712 555620 234764 555626
rect 234712 555562 234764 555568
rect 234908 555558 234936 556430
rect 235828 556102 235856 559098
rect 235908 559020 235960 559026
rect 235908 558962 235960 558968
rect 235920 556102 235948 558962
rect 237392 556594 237420 630634
rect 255332 576854 255360 700402
rect 267660 700398 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 256700 700392 256752 700398
rect 256700 700334 256752 700340
rect 267648 700392 267700 700398
rect 267648 700334 267700 700340
rect 256712 576854 256740 700334
rect 255332 576826 255912 576854
rect 256712 576826 257200 576854
rect 238760 562148 238812 562154
rect 238760 562090 238812 562096
rect 238772 556594 238800 562090
rect 253296 562080 253348 562086
rect 253296 562022 253348 562028
rect 241704 561740 241756 561746
rect 241704 561682 241756 561688
rect 241152 557728 241204 557734
rect 241152 557670 241204 557676
rect 241164 556594 241192 557670
rect 237392 556566 237636 556594
rect 238772 556566 238924 556594
rect 240856 556566 241192 556594
rect 241716 556594 241744 561682
rect 252008 560992 252060 560998
rect 252008 560934 252060 560940
rect 244280 560448 244332 560454
rect 244280 560390 244332 560396
rect 243404 556608 243460 556617
rect 241716 556566 242144 556594
rect 244292 556594 244320 560390
rect 249800 560380 249852 560386
rect 249800 560322 249852 560328
rect 245660 559700 245712 559706
rect 245660 559642 245712 559648
rect 245672 556594 245700 559642
rect 248558 556776 248610 556782
rect 248558 556718 248610 556724
rect 244292 556566 244720 556594
rect 245672 556566 246008 556594
rect 248570 556580 248598 556718
rect 249812 556594 249840 560322
rect 251086 557560 251142 557569
rect 251086 557495 251142 557504
rect 251100 556594 251128 557495
rect 252020 556594 252048 560934
rect 253308 556594 253336 562022
rect 255884 556594 255912 576826
rect 257172 556594 257200 576826
rect 282932 570722 282960 702406
rect 300136 699718 300164 703520
rect 332520 700466 332548 703520
rect 348804 702434 348832 703520
rect 364996 702434 365024 703520
rect 347792 702406 348832 702434
rect 364352 702406 365024 702434
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 306380 699712 306432 699718
rect 306380 699654 306432 699660
rect 298100 670812 298152 670818
rect 298100 670754 298152 670760
rect 293960 616888 294012 616894
rect 293960 616830 294012 616836
rect 293972 576854 294000 616830
rect 293972 576826 294552 576854
rect 282920 570716 282972 570722
rect 282920 570658 282972 570664
rect 260380 562012 260432 562018
rect 260380 561954 260432 561960
rect 259460 557796 259512 557802
rect 259460 557738 259512 557744
rect 259472 556594 259500 557738
rect 260392 556594 260420 561954
rect 279056 561944 279108 561950
rect 279056 561886 279108 561892
rect 270684 561876 270736 561882
rect 270684 561818 270736 561824
rect 273260 561876 273312 561882
rect 273260 561818 273312 561824
rect 268108 560652 268160 560658
rect 268108 560594 268160 560600
rect 261668 559700 261720 559706
rect 261668 559642 261720 559648
rect 249812 556566 249872 556594
rect 251100 556566 251160 556594
rect 252020 556566 252448 556594
rect 253308 556566 253736 556594
rect 255884 556566 256312 556594
rect 257172 556566 257600 556594
rect 259472 556566 259532 556594
rect 260392 556566 260820 556594
rect 243404 556543 243460 556552
rect 247052 556306 247296 556322
rect 247040 556300 247296 556306
rect 247092 556294 247296 556300
rect 247040 556242 247092 556248
rect 254676 556232 254728 556238
rect 254728 556180 255024 556186
rect 254676 556174 255024 556180
rect 254688 556158 255024 556174
rect 261680 556102 261708 559642
rect 263048 559496 263100 559502
rect 263048 559438 263100 559444
rect 261760 559020 261812 559026
rect 261760 558962 261812 558968
rect 262864 559020 262916 559026
rect 262864 558962 262916 558968
rect 261772 556594 261800 558962
rect 262876 558278 262904 558962
rect 262864 558272 262916 558278
rect 262864 558214 262916 558220
rect 263060 556594 263088 559438
rect 265624 558952 265676 558958
rect 265624 558894 265676 558900
rect 265636 556594 265664 558894
rect 266912 556980 266964 556986
rect 266912 556922 266964 556928
rect 266924 556594 266952 556922
rect 268120 556594 268148 560594
rect 269488 556640 269540 556646
rect 261772 556566 262108 556594
rect 263060 556566 263396 556594
rect 265636 556566 265972 556594
rect 266924 556566 267260 556594
rect 268120 556566 268548 556594
rect 270696 556594 270724 561818
rect 271972 560788 272024 560794
rect 271972 560730 272024 560736
rect 271984 556594 272012 560730
rect 273272 556594 273300 561818
rect 274732 559496 274784 559502
rect 274732 559438 274784 559444
rect 274640 559020 274692 559026
rect 274640 558962 274692 558968
rect 274652 556594 274680 558962
rect 274744 558346 274772 559438
rect 274732 558340 274784 558346
rect 274732 558282 274784 558288
rect 277858 557832 277914 557841
rect 277858 557767 277914 557776
rect 277872 556594 277900 557767
rect 269540 556588 269836 556594
rect 269488 556582 269836 556588
rect 269500 556566 269836 556582
rect 270696 556566 271124 556594
rect 271984 556566 272412 556594
rect 273272 556566 273700 556594
rect 274652 556566 274988 556594
rect 277564 556566 277900 556594
rect 279068 556594 279096 561886
rect 293224 560788 293276 560794
rect 293224 560730 293276 560736
rect 280344 560584 280396 560590
rect 280344 560526 280396 560532
rect 280356 556594 280384 560526
rect 289452 559632 289504 559638
rect 289452 559574 289504 559580
rect 288440 559564 288492 559570
rect 288440 559506 288492 559512
rect 284300 558476 284352 558482
rect 284300 558418 284352 558424
rect 282044 556880 282100 556889
rect 282044 556815 282100 556824
rect 279068 556566 279496 556594
rect 280356 556566 280784 556594
rect 282058 556580 282086 556815
rect 284312 556594 284340 558418
rect 287060 558408 287112 558414
rect 287060 558350 287112 558356
rect 285680 557864 285732 557870
rect 285680 557806 285732 557812
rect 285692 556594 285720 557806
rect 287072 556594 287100 558350
rect 288452 556594 288480 559506
rect 289464 556594 289492 559574
rect 292028 559360 292080 559366
rect 292028 559302 292080 559308
rect 292040 556594 292068 559302
rect 293236 556594 293264 560730
rect 294524 556594 294552 576826
rect 298112 556594 298140 670754
rect 306392 576854 306420 699654
rect 340880 683188 340932 683194
rect 340880 683130 340932 683136
rect 314660 618316 314712 618322
rect 314660 618258 314712 618264
rect 306392 576826 306788 576854
rect 305460 574796 305512 574802
rect 305460 574738 305512 574744
rect 302884 560652 302936 560658
rect 302884 560594 302936 560600
rect 300308 560584 300360 560590
rect 300308 560526 300360 560532
rect 299432 556880 299488 556889
rect 299432 556815 299488 556824
rect 284312 556566 284648 556594
rect 285692 556566 285936 556594
rect 287072 556566 287224 556594
rect 288452 556566 288512 556594
rect 289464 556566 289800 556594
rect 292040 556566 292376 556594
rect 293236 556566 293664 556594
rect 294524 556566 294952 556594
rect 298112 556566 298172 556594
rect 299446 556580 299474 556815
rect 300320 556594 300348 560526
rect 301688 559700 301740 559706
rect 301688 559642 301740 559648
rect 301700 556594 301728 559642
rect 302896 556594 302924 560594
rect 304906 559328 304962 559337
rect 304906 559263 304962 559272
rect 304920 556594 304948 559263
rect 300320 556566 300748 556594
rect 301700 556566 302036 556594
rect 302896 556566 303324 556594
rect 304612 556566 304948 556594
rect 305472 556594 305500 574738
rect 306760 556594 306788 576826
rect 309324 560856 309376 560862
rect 309324 560798 309376 560804
rect 308772 557796 308824 557802
rect 308772 557738 308824 557744
rect 308784 556594 308812 557738
rect 305472 556566 305900 556594
rect 306760 556566 307188 556594
rect 308476 556566 308812 556594
rect 309336 556594 309364 560798
rect 312636 556640 312688 556646
rect 309336 556566 309764 556594
rect 312340 556588 312636 556594
rect 312340 556582 312688 556588
rect 314672 556594 314700 618258
rect 340892 576854 340920 683130
rect 340892 576826 341564 576854
rect 340236 562216 340288 562222
rect 340236 562158 340288 562164
rect 324320 561808 324372 561814
rect 324320 561750 324372 561756
rect 316040 560924 316092 560930
rect 316040 560866 316092 560872
rect 316052 556594 316080 560866
rect 322940 559428 322992 559434
rect 322940 559370 322992 559376
rect 320364 558136 320416 558142
rect 320364 558078 320416 558084
rect 317788 557932 317840 557938
rect 317788 557874 317840 557880
rect 317800 556594 317828 557874
rect 320376 556594 320404 558078
rect 321652 556708 321704 556714
rect 321652 556650 321704 556656
rect 321664 556594 321692 556650
rect 322952 556594 322980 559370
rect 324332 556594 324360 561750
rect 329288 560924 329340 560930
rect 329288 560866 329340 560872
rect 328092 558068 328144 558074
rect 328092 558010 328144 558016
rect 327078 557152 327134 557161
rect 327078 557087 327134 557096
rect 327092 556594 327120 557087
rect 328104 556594 328132 558010
rect 329300 556594 329328 560866
rect 334440 560516 334492 560522
rect 334440 560458 334492 560464
rect 330666 558104 330722 558113
rect 330666 558039 330722 558048
rect 330680 556594 330708 558039
rect 333566 556776 333618 556782
rect 333566 556718 333618 556724
rect 332508 556708 332560 556714
rect 332508 556650 332560 556656
rect 332520 556594 332548 556650
rect 312340 556566 312676 556582
rect 314672 556566 314916 556594
rect 316052 556566 316204 556594
rect 317800 556566 318136 556594
rect 320376 556566 320712 556594
rect 321664 556566 322000 556594
rect 322952 556566 323288 556594
rect 324332 556566 324576 556594
rect 327092 556566 327152 556594
rect 328104 556566 328440 556594
rect 329300 556566 329728 556594
rect 330680 556566 331016 556594
rect 332304 556566 332548 556594
rect 333578 556580 333606 556718
rect 334452 556594 334480 560458
rect 340248 556594 340276 562158
rect 341536 556594 341564 576826
rect 345388 565888 345440 565894
rect 345388 565830 345440 565836
rect 343548 558272 343600 558278
rect 343548 558214 343600 558220
rect 343560 556594 343588 558214
rect 344836 557932 344888 557938
rect 344836 557874 344888 557880
rect 344848 556594 344876 557874
rect 334452 556566 334880 556594
rect 339388 556578 339540 556594
rect 339388 556572 339552 556578
rect 339388 556566 339500 556572
rect 340248 556566 340676 556594
rect 341536 556566 341964 556594
rect 343252 556566 343588 556594
rect 344540 556566 344876 556594
rect 345400 556594 345428 565830
rect 347792 563786 347820 702406
rect 347780 563780 347832 563786
rect 347780 563722 347832 563728
rect 364352 563718 364380 702406
rect 397472 700534 397500 703520
rect 397460 700528 397512 700534
rect 397460 700470 397512 700476
rect 407120 700460 407172 700466
rect 407120 700402 407172 700408
rect 407132 576854 407160 700402
rect 407132 576826 407896 576854
rect 364340 563712 364392 563718
rect 364340 563654 364392 563660
rect 406568 563100 406620 563106
rect 406568 563042 406620 563048
rect 371792 562556 371844 562562
rect 371792 562498 371844 562504
rect 350540 561060 350592 561066
rect 350540 561002 350592 561008
rect 347962 560552 348018 560561
rect 347962 560487 348018 560496
rect 346766 559872 346822 559881
rect 346766 559807 346822 559816
rect 346780 556594 346808 559807
rect 347976 556594 348004 560487
rect 349988 558136 350040 558142
rect 349988 558078 350040 558084
rect 350000 556594 350028 558078
rect 345400 556566 345828 556594
rect 346780 556566 347116 556594
rect 347976 556566 348404 556594
rect 349692 556566 350028 556594
rect 350552 556594 350580 561002
rect 360936 559972 360988 559978
rect 360936 559914 360988 559920
rect 358358 559872 358414 559881
rect 358358 559807 358414 559816
rect 354680 559292 354732 559298
rect 354680 559234 354732 559240
rect 353300 557184 353352 557190
rect 353300 557126 353352 557132
rect 353312 556594 353340 557126
rect 354692 556594 354720 559234
rect 356428 558000 356480 558006
rect 356428 557942 356480 557948
rect 356440 556594 356468 557942
rect 358372 556594 358400 559807
rect 360948 556850 360976 559914
rect 368020 559904 368072 559910
rect 368020 559846 368072 559852
rect 365810 559736 365866 559745
rect 365810 559671 365866 559680
rect 362960 559496 363012 559502
rect 362960 559438 363012 559444
rect 360936 556844 360988 556850
rect 360936 556786 360988 556792
rect 350552 556566 350980 556594
rect 353312 556566 353556 556594
rect 354692 556566 354844 556594
rect 356440 556566 356776 556594
rect 358064 556566 358400 556594
rect 362972 556594 363000 559438
rect 365824 556730 365852 559671
rect 367008 559224 367060 559230
rect 367008 559166 367060 559172
rect 367020 558249 367048 559166
rect 367006 558240 367062 558249
rect 367006 558175 367062 558184
rect 366732 557048 366784 557054
rect 366732 556990 366784 556996
rect 365778 556702 365852 556730
rect 362972 556566 363216 556594
rect 365778 556580 365806 556702
rect 366744 556594 366772 556990
rect 368032 556594 368060 559846
rect 369308 557116 369360 557122
rect 369308 557058 369360 557064
rect 369320 556594 369348 557058
rect 370918 556844 370970 556850
rect 370918 556786 370970 556792
rect 366744 556566 367080 556594
rect 368032 556566 368368 556594
rect 369320 556566 369656 556594
rect 370930 556580 370958 556786
rect 371804 556594 371832 562498
rect 382740 560720 382792 560726
rect 382740 560662 382792 560668
rect 375378 559600 375434 559609
rect 375378 559535 375434 559544
rect 373170 557016 373226 557025
rect 373170 556951 373226 556960
rect 373184 556594 373212 556951
rect 375392 556594 375420 559535
rect 378968 559156 379020 559162
rect 378968 559098 379020 559104
rect 377680 559088 377732 559094
rect 377680 559030 377732 559036
rect 378784 559088 378836 559094
rect 378784 559030 378836 559036
rect 376668 557048 376720 557054
rect 376668 556990 376720 556996
rect 376680 556594 376708 556990
rect 377692 556594 377720 559030
rect 378796 558210 378824 559030
rect 378784 558204 378836 558210
rect 378784 558146 378836 558152
rect 378980 556594 379008 559098
rect 382752 556594 382780 560662
rect 388628 559904 388680 559910
rect 388628 559846 388680 559852
rect 384118 559464 384174 559473
rect 384118 559399 384174 559408
rect 384132 556594 384160 559399
rect 386052 557116 386104 557122
rect 386052 557058 386104 557064
rect 386064 556594 386092 557058
rect 387340 556980 387392 556986
rect 387340 556922 387392 556928
rect 387352 556594 387380 556922
rect 388640 556594 388668 559846
rect 393412 559836 393464 559842
rect 393412 559778 393464 559784
rect 389272 559224 389324 559230
rect 389272 559166 389324 559172
rect 371804 556566 372232 556594
rect 373184 556566 373520 556594
rect 375392 556566 375452 556594
rect 376680 556566 376740 556594
rect 377692 556566 378028 556594
rect 378980 556566 379316 556594
rect 382752 556566 383180 556594
rect 384132 556566 384468 556594
rect 385756 556566 386092 556594
rect 387044 556566 387380 556594
rect 388332 556566 388668 556594
rect 389284 556594 389312 559166
rect 392492 559156 392544 559162
rect 392492 559098 392544 559104
rect 391204 557864 391256 557870
rect 391204 557806 391256 557812
rect 391216 556594 391244 557806
rect 392504 556594 392532 559098
rect 393320 558952 393372 558958
rect 393320 558894 393372 558900
rect 393332 556918 393360 558894
rect 393320 556912 393372 556918
rect 393320 556854 393372 556860
rect 389284 556566 389620 556594
rect 390908 556566 391244 556594
rect 392196 556566 392532 556594
rect 393424 556594 393452 559778
rect 402152 559360 402204 559366
rect 402152 559302 402204 559308
rect 398288 559020 398340 559026
rect 398288 558962 398340 558968
rect 398300 556594 398328 558962
rect 400864 558204 400916 558210
rect 400864 558146 400916 558152
rect 400876 556594 400904 558146
rect 402164 556594 402192 559302
rect 403440 559224 403492 559230
rect 403440 559166 403492 559172
rect 403452 556594 403480 559166
rect 404728 558000 404780 558006
rect 404728 557942 404780 557948
rect 404740 556594 404768 557942
rect 405372 557592 405424 557598
rect 405372 557534 405424 557540
rect 393424 556566 393484 556594
rect 397992 556566 398328 556594
rect 400568 556566 400904 556594
rect 401856 556566 402192 556594
rect 403144 556566 403480 556594
rect 404432 556566 404768 556594
rect 405384 556594 405412 557534
rect 406580 556594 406608 563042
rect 407868 556594 407896 576826
rect 412652 572014 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429212 574802 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 459652 700528 459704 700534
rect 459652 700470 459704 700476
rect 436100 700392 436152 700398
rect 436100 700334 436152 700340
rect 436112 576854 436140 700334
rect 452660 670744 452712 670750
rect 452660 670686 452712 670692
rect 436112 576826 436232 576854
rect 429200 574796 429252 574802
rect 429200 574738 429252 574744
rect 412640 572008 412692 572014
rect 412640 571950 412692 571956
rect 426532 562488 426584 562494
rect 426532 562430 426584 562436
rect 414938 560416 414994 560425
rect 414938 560351 414994 560360
rect 414388 559564 414440 559570
rect 414388 559506 414440 559512
rect 412456 559496 412508 559502
rect 412456 559438 412508 559444
rect 409234 559056 409290 559065
rect 409234 558991 409290 559000
rect 409248 556594 409276 558991
rect 410522 557968 410578 557977
rect 410522 557903 410578 557912
rect 410536 556594 410564 557903
rect 412468 556594 412496 559438
rect 414400 556594 414428 559506
rect 405384 556566 405720 556594
rect 406580 556566 407008 556594
rect 407868 556566 408296 556594
rect 409248 556566 409584 556594
rect 410536 556566 410872 556594
rect 412160 556566 412496 556594
rect 414092 556566 414428 556594
rect 414952 556594 414980 560351
rect 424048 559768 424100 559774
rect 424048 559710 424100 559716
rect 419448 559700 419500 559706
rect 419448 559642 419500 559648
rect 416688 559632 416740 559638
rect 416688 559574 416740 559580
rect 416700 556730 416728 559574
rect 417606 559192 417662 559201
rect 417606 559127 417662 559136
rect 416654 556702 416728 556730
rect 414952 556566 415380 556594
rect 416654 556580 416682 556702
rect 417620 556594 417648 559127
rect 419460 556594 419488 559642
rect 420828 559428 420880 559434
rect 420828 559370 420880 559376
rect 420840 556594 420868 559370
rect 421472 558952 421524 558958
rect 421472 558894 421524 558900
rect 423404 558952 423456 558958
rect 423404 558894 423456 558900
rect 417620 556566 417956 556594
rect 419244 556566 419488 556594
rect 420532 556566 420868 556594
rect 421484 556594 421512 558894
rect 423416 556594 423444 558894
rect 421484 556566 421820 556594
rect 423108 556566 423444 556594
rect 424060 556594 424088 559710
rect 425980 556912 426032 556918
rect 425980 556854 426032 556860
rect 425992 556594 426020 556854
rect 424060 556566 424396 556594
rect 425684 556566 426020 556594
rect 426544 556594 426572 562430
rect 430580 559088 430632 559094
rect 430580 559030 430632 559036
rect 432420 559088 432472 559094
rect 432420 559030 432472 559036
rect 429198 557696 429254 557705
rect 429198 557631 429254 557640
rect 429212 556594 429240 557631
rect 430592 556594 430620 559030
rect 432432 556594 432460 559030
rect 433708 557660 433760 557666
rect 433708 557602 433760 557608
rect 426544 556566 426972 556594
rect 429212 556566 429548 556594
rect 430592 556566 430836 556594
rect 432124 556566 432460 556594
rect 433720 556594 433748 557602
rect 435640 557592 435692 557598
rect 435640 557534 435692 557540
rect 435652 556594 435680 557534
rect 433720 556566 434056 556594
rect 435344 556566 435680 556594
rect 436204 556594 436232 576826
rect 441620 562284 441672 562290
rect 441620 562226 441672 562232
rect 440790 559600 440846 559609
rect 440790 559535 440846 559544
rect 438216 559292 438268 559298
rect 438216 559234 438268 559240
rect 438228 556594 438256 559234
rect 439502 559192 439558 559201
rect 439502 559127 439558 559136
rect 439516 556594 439544 559127
rect 440804 556594 440832 559535
rect 436204 556566 436632 556594
rect 437920 556566 438256 556594
rect 439208 556566 439544 556594
rect 440496 556566 440832 556594
rect 441632 556594 441660 562226
rect 445208 560312 445260 560318
rect 445208 560254 445260 560260
rect 444286 559464 444342 559473
rect 444286 559399 444342 559408
rect 443368 557660 443420 557666
rect 443368 557602 443420 557608
rect 443380 556594 443408 557602
rect 441632 556566 441784 556594
rect 443072 556566 443408 556594
rect 444300 556594 444328 559399
rect 445220 556594 445248 560254
rect 446588 559972 446640 559978
rect 446588 559914 446640 559920
rect 446600 556594 446628 559914
rect 451740 559904 451792 559910
rect 451740 559846 451792 559852
rect 451648 559156 451700 559162
rect 451648 559098 451700 559104
rect 448426 559056 448482 559065
rect 448426 558991 448482 559000
rect 448440 556594 448468 558991
rect 449808 558068 449860 558074
rect 449808 558010 449860 558016
rect 449820 556594 449848 558010
rect 451556 557048 451608 557054
rect 451556 556990 451608 556996
rect 450772 556744 450828 556753
rect 450772 556679 450828 556688
rect 444300 556566 444360 556594
rect 445220 556566 445648 556594
rect 446600 556566 446936 556594
rect 448224 556566 448468 556594
rect 449512 556566 449848 556594
rect 450786 556580 450814 556679
rect 339500 556514 339552 556520
rect 359004 556504 359056 556510
rect 313600 556472 313656 556481
rect 283024 556442 283360 556458
rect 283012 556436 283360 556442
rect 283064 556430 283360 556436
rect 291088 556442 291240 556458
rect 291088 556436 291252 556442
rect 291088 556430 291200 556436
rect 283012 556378 283064 556384
rect 313600 556407 313656 556416
rect 319396 556472 319452 556481
rect 360936 556504 360988 556510
rect 359056 556452 359352 556458
rect 359004 556446 359352 556452
rect 359016 556430 359352 556446
rect 360640 556452 360936 556458
rect 360640 556446 360988 556452
rect 360640 556430 360976 556446
rect 319396 556407 319452 556416
rect 291200 556378 291252 556384
rect 276020 556368 276072 556374
rect 296444 556368 296496 556374
rect 276072 556316 276276 556322
rect 276020 556310 276276 556316
rect 276032 556294 276276 556310
rect 296240 556316 296444 556322
rect 296240 556310 296496 556316
rect 325836 556336 325892 556345
rect 296240 556294 296484 556310
rect 395416 556306 395752 556322
rect 395416 556300 395764 556306
rect 395416 556294 395712 556300
rect 325836 556271 325892 556280
rect 395712 556242 395764 556248
rect 399576 556232 399628 556238
rect 399280 556180 399576 556186
rect 399280 556174 399628 556180
rect 399280 556158 399616 556174
rect 235816 556096 235868 556102
rect 235032 556064 235088 556073
rect 235816 556038 235868 556044
rect 235908 556096 235960 556102
rect 235908 556038 235960 556044
rect 261668 556096 261720 556102
rect 364800 556096 364852 556102
rect 261668 556038 261720 556044
rect 364504 556044 364800 556050
rect 364504 556038 364852 556044
rect 364504 556022 364840 556038
rect 235032 555999 235088 556008
rect 236320 555928 236376 555937
rect 236320 555863 236376 555872
rect 264656 555928 264712 555937
rect 264656 555863 264712 555872
rect 338072 555928 338128 555937
rect 338072 555863 338128 555872
rect 352240 555928 352296 555937
rect 352240 555863 352296 555872
rect 234896 555552 234948 555558
rect 234896 555494 234948 555500
rect 234710 417616 234766 417625
rect 234710 417551 234766 417560
rect 234620 395344 234672 395350
rect 234620 395286 234672 395292
rect 234724 335354 234752 417551
rect 234802 370016 234858 370025
rect 234802 369951 234858 369960
rect 234632 335326 234752 335354
rect 234632 334762 234660 335326
rect 234620 334756 234672 334762
rect 234620 334698 234672 334704
rect 234816 332042 234844 369951
rect 236000 338224 236052 338230
rect 447140 338224 447192 338230
rect 236000 338166 236052 338172
rect 240506 338192 240562 338201
rect 234908 338014 235060 338042
rect 234908 335918 234936 338014
rect 234896 335912 234948 335918
rect 234896 335854 234948 335860
rect 234804 332036 234856 332042
rect 234804 331978 234856 331984
rect 234528 273216 234580 273222
rect 234528 273158 234580 273164
rect 234620 47592 234672 47598
rect 234620 47534 234672 47540
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 480 234660 47534
rect 235816 13116 235868 13122
rect 235816 13058 235868 13064
rect 235828 480 235856 13058
rect 236012 490 236040 338166
rect 240506 338127 240562 338136
rect 267738 338192 267794 338201
rect 267738 338127 267794 338136
rect 270774 338192 270830 338201
rect 270774 338127 270830 338136
rect 379518 338192 379574 338201
rect 379518 338127 379574 338136
rect 398930 338192 398986 338201
rect 412362 338192 412418 338201
rect 412160 338150 412362 338178
rect 398930 338127 398986 338136
rect 447140 338166 447192 338172
rect 450358 338192 450414 338201
rect 412362 338127 412418 338136
rect 236104 338014 236348 338042
rect 237484 338014 237636 338042
rect 238864 338014 238924 338042
rect 236104 4962 236132 338014
rect 237378 337920 237434 337929
rect 237378 337855 237434 337864
rect 237392 16574 237420 337855
rect 237484 32434 237512 338014
rect 238758 337648 238814 337657
rect 238758 337583 238814 337592
rect 237472 32428 237524 32434
rect 237472 32370 237524 32376
rect 237392 16546 237696 16574
rect 236092 4956 236144 4962
rect 236092 4898 236144 4904
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236012 462 236592 490
rect 236564 354 236592 462
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 238772 3482 238800 337583
rect 238864 5166 238892 338014
rect 240198 337770 240226 338028
rect 240198 337742 240272 337770
rect 238852 5160 238904 5166
rect 238852 5102 238904 5108
rect 240244 4894 240272 337742
rect 240520 335354 240548 338127
rect 241164 338014 241500 338042
rect 242360 338014 242788 338042
rect 243004 338014 244076 338042
rect 245028 338014 245364 338042
rect 246316 338014 246652 338042
rect 247512 338014 247940 338042
rect 248800 338014 249228 338042
rect 250088 338014 250516 338042
rect 251376 338014 251804 338042
rect 253092 338014 253428 338042
rect 255024 338014 255268 338042
rect 241164 336598 241192 338014
rect 241152 336592 241204 336598
rect 241152 336534 241204 336540
rect 240336 335326 240548 335354
rect 240232 4888 240284 4894
rect 240232 4830 240284 4836
rect 238772 3454 239352 3482
rect 239324 480 239352 3454
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240336 354 240364 335326
rect 241520 334756 241572 334762
rect 241520 334698 241572 334704
rect 241532 16574 241560 334698
rect 242360 316034 242388 338014
rect 241624 316006 242388 316034
rect 241624 57254 241652 316006
rect 243004 290562 243032 338014
rect 244280 337680 244332 337686
rect 244280 337622 244332 337628
rect 243084 337408 243136 337414
rect 243084 337350 243136 337356
rect 242992 290556 243044 290562
rect 242992 290498 243044 290504
rect 241612 57248 241664 57254
rect 241612 57190 241664 57196
rect 243096 16574 243124 337350
rect 244292 16574 244320 337622
rect 245028 336870 245056 338014
rect 245016 336864 245068 336870
rect 245016 336806 245068 336812
rect 246316 336598 246344 338014
rect 244924 336592 244976 336598
rect 244924 336534 244976 336540
rect 246304 336592 246356 336598
rect 246304 336534 246356 336540
rect 244936 158030 244964 336534
rect 247512 316034 247540 338014
rect 248420 333464 248472 333470
rect 248420 333406 248472 333412
rect 247052 316006 247540 316034
rect 247052 179382 247080 316006
rect 247040 179376 247092 179382
rect 247040 179318 247092 179324
rect 244924 158024 244976 158030
rect 244924 157966 244976 157972
rect 241532 16546 241744 16574
rect 243096 16546 244136 16574
rect 244292 16546 245240 16574
rect 241716 480 241744 16546
rect 242900 3256 242952 3262
rect 242900 3198 242952 3204
rect 242912 480 242940 3198
rect 244108 480 244136 16546
rect 245212 480 245240 16546
rect 247592 6724 247644 6730
rect 247592 6666 247644 6672
rect 246396 3324 246448 3330
rect 246396 3266 246448 3272
rect 246408 480 246436 3266
rect 247604 480 247632 6666
rect 240478 354 240590 480
rect 240336 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 333406
rect 248800 316034 248828 338014
rect 249800 337408 249852 337414
rect 249800 337350 249852 337356
rect 248524 316006 248828 316034
rect 248524 5030 248552 316006
rect 248512 5024 248564 5030
rect 248512 4966 248564 4972
rect 249812 3482 249840 337350
rect 250088 316034 250116 338014
rect 251180 326460 251232 326466
rect 251180 326402 251232 326408
rect 249904 316006 250116 316034
rect 249904 3738 249932 316006
rect 249892 3732 249944 3738
rect 249892 3674 249944 3680
rect 249812 3454 250024 3482
rect 249996 480 250024 3454
rect 251192 480 251220 326402
rect 251376 316034 251404 338014
rect 253400 333674 253428 338014
rect 253940 337612 253992 337618
rect 253940 337554 253992 337560
rect 253388 333668 253440 333674
rect 253388 333610 253440 333616
rect 251284 316006 251404 316034
rect 251284 291854 251312 316006
rect 251272 291848 251324 291854
rect 251272 291790 251324 291796
rect 253952 16574 253980 337554
rect 255240 333742 255268 338014
rect 255884 338014 256312 338042
rect 257172 338014 257600 338042
rect 258460 338014 258888 338042
rect 259564 338014 260176 338042
rect 262416 338014 262752 338042
rect 263612 338014 264040 338042
rect 264992 338014 265328 338042
rect 266372 338014 266616 338042
rect 255228 333736 255280 333742
rect 255228 333678 255280 333684
rect 255884 316034 255912 338014
rect 257172 316034 257200 338014
rect 258460 316034 258488 338014
rect 255332 316006 255912 316034
rect 256712 316006 257200 316034
rect 258092 316006 258488 316034
rect 255332 272542 255360 316006
rect 255320 272536 255372 272542
rect 255320 272478 255372 272484
rect 253952 16546 254256 16574
rect 252376 5976 252428 5982
rect 252376 5918 252428 5924
rect 252388 480 252416 5918
rect 253480 4888 253532 4894
rect 253480 4830 253532 4836
rect 253492 480 253520 4830
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255872 6316 255924 6322
rect 255872 6258 255924 6264
rect 255884 480 255912 6258
rect 256712 5982 256740 316006
rect 256700 5976 256752 5982
rect 256700 5918 256752 5924
rect 258092 5098 258120 316006
rect 259564 300218 259592 338014
rect 262220 337544 262272 337550
rect 262220 337486 262272 337492
rect 259644 334756 259696 334762
rect 259644 334698 259696 334704
rect 259552 300212 259604 300218
rect 259552 300154 259604 300160
rect 259656 6914 259684 334698
rect 260840 315376 260892 315382
rect 260840 315318 260892 315324
rect 260852 16574 260880 315318
rect 262232 16574 262260 337486
rect 262416 336802 262444 338014
rect 262404 336796 262456 336802
rect 262404 336738 262456 336744
rect 263612 123486 263640 338014
rect 263600 123480 263652 123486
rect 263600 123422 263652 123428
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 259472 6886 259684 6914
rect 258264 6316 258316 6322
rect 258264 6258 258316 6264
rect 258080 5092 258132 5098
rect 258080 5034 258132 5040
rect 257068 5024 257120 5030
rect 257068 4966 257120 4972
rect 257080 480 257108 4966
rect 258276 480 258304 6258
rect 259472 480 259500 6886
rect 260656 3392 260708 3398
rect 260656 3334 260708 3340
rect 260668 480 260696 3334
rect 261772 480 261800 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264992 9042 265020 338014
rect 266372 336666 266400 338014
rect 266360 336660 266412 336666
rect 266360 336602 266412 336608
rect 266358 327856 266414 327865
rect 266358 327791 266414 327800
rect 266372 16574 266400 327791
rect 266372 16546 266584 16574
rect 264980 9036 265032 9042
rect 264980 8978 265032 8984
rect 264152 4140 264204 4146
rect 264152 4082 264204 4088
rect 264164 480 264192 4082
rect 265348 3732 265400 3738
rect 265348 3674 265400 3680
rect 265360 480 265388 3674
rect 266556 480 266584 16546
rect 267752 480 267780 338127
rect 267890 337770 267918 338028
rect 269132 338014 269192 338042
rect 270052 338014 270480 338042
rect 267890 337742 267964 337770
rect 267832 331900 267884 331906
rect 267832 331842 267884 331848
rect 267844 16574 267872 331842
rect 267936 97986 267964 337742
rect 269132 336326 269160 338014
rect 269120 336320 269172 336326
rect 269120 336262 269172 336268
rect 270052 316034 270080 338014
rect 270788 335354 270816 338127
rect 270696 335326 270816 335354
rect 271432 338014 271768 338042
rect 273272 338014 273700 338042
rect 274988 338014 275324 338042
rect 270592 330472 270644 330478
rect 270592 330414 270644 330420
rect 269316 316006 270080 316034
rect 267924 97980 267976 97986
rect 267924 97922 267976 97928
rect 269316 51814 269344 316006
rect 269304 51808 269356 51814
rect 269304 51750 269356 51756
rect 269212 51740 269264 51746
rect 269212 51682 269264 51688
rect 269224 16574 269252 51682
rect 267844 16546 268424 16574
rect 269224 16546 270080 16574
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 270604 11762 270632 330414
rect 270696 16574 270724 335326
rect 271432 330478 271460 338014
rect 271880 332036 271932 332042
rect 271880 331978 271932 331984
rect 271420 330472 271472 330478
rect 271420 330414 271472 330420
rect 271892 16574 271920 331978
rect 270696 16546 270816 16574
rect 271892 16546 272472 16574
rect 270592 11756 270644 11762
rect 270592 11698 270644 11704
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 273272 8022 273300 338014
rect 275296 333606 275324 338014
rect 276124 338014 276276 338042
rect 277504 338014 277564 338042
rect 279712 338014 280140 338042
rect 280724 338014 281428 338042
rect 282380 338014 282716 338042
rect 283668 338014 284004 338042
rect 284864 338014 285292 338042
rect 286580 338014 286916 338042
rect 275376 336592 275428 336598
rect 275376 336534 275428 336540
rect 275284 333600 275336 333606
rect 275284 333542 275336 333548
rect 275388 316034 275416 336534
rect 276020 318096 276072 318102
rect 276020 318038 276072 318044
rect 275296 316006 275416 316034
rect 275296 145586 275324 316006
rect 275284 145580 275336 145586
rect 275284 145522 275336 145528
rect 276032 16574 276060 318038
rect 276124 29646 276152 338014
rect 277400 336320 277452 336326
rect 277400 336262 277452 336268
rect 276112 29640 276164 29646
rect 276112 29582 276164 29588
rect 276032 16546 276704 16574
rect 273352 13184 273404 13190
rect 273352 13126 273404 13132
rect 273260 8016 273312 8022
rect 273260 7958 273312 7964
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273364 354 273392 13126
rect 276020 6044 276072 6050
rect 276020 5986 276072 5992
rect 274824 5160 274876 5166
rect 274824 5102 274876 5108
rect 274836 480 274864 5102
rect 276032 480 276060 5986
rect 273598 354 273710 480
rect 273364 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 277412 6914 277440 336262
rect 277504 7682 277532 338014
rect 278780 337476 278832 337482
rect 278780 337418 278832 337424
rect 278792 16574 278820 337418
rect 279712 316034 279740 338014
rect 280160 323604 280212 323610
rect 280160 323546 280212 323552
rect 278884 316006 279740 316034
rect 278884 232558 278912 316006
rect 278872 232552 278924 232558
rect 278872 232494 278924 232500
rect 280172 16574 280200 323546
rect 280724 316034 280752 338014
rect 282380 335986 282408 338014
rect 283668 336598 283696 338014
rect 283656 336592 283708 336598
rect 283656 336534 283708 336540
rect 280804 335980 280856 335986
rect 280804 335922 280856 335928
rect 282368 335980 282420 335986
rect 282368 335922 282420 335928
rect 280264 316006 280752 316034
rect 280264 280838 280292 316006
rect 280252 280832 280304 280838
rect 280252 280774 280304 280780
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 277492 7676 277544 7682
rect 277492 7618 277544 7624
rect 277412 6886 278360 6914
rect 278332 480 278360 6886
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 280816 3602 280844 335922
rect 282920 334960 282972 334966
rect 282920 334902 282972 334908
rect 281540 330608 281592 330614
rect 281540 330550 281592 330556
rect 280804 3596 280856 3602
rect 280804 3538 280856 3544
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 330550
rect 282932 16574 282960 334902
rect 284300 327820 284352 327826
rect 284300 327762 284352 327768
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 480 284340 327762
rect 284392 318096 284444 318102
rect 284392 318038 284444 318044
rect 284404 16574 284432 318038
rect 284864 316034 284892 338014
rect 286888 333878 286916 338014
rect 287440 338014 287868 338042
rect 288728 338014 289156 338042
rect 291304 338014 291732 338042
rect 293236 338014 293664 338042
rect 294524 338014 294952 338042
rect 295812 338014 296240 338042
rect 297100 338014 297528 338042
rect 298388 338014 298816 338042
rect 299676 338014 300104 338042
rect 300964 338014 301392 338042
rect 302344 338014 302680 338042
rect 305012 338014 305256 338042
rect 306392 338014 306544 338042
rect 286876 333872 286928 333878
rect 286876 333814 286928 333820
rect 287440 316034 287468 338014
rect 288728 316034 288756 338014
rect 291200 336524 291252 336530
rect 291200 336466 291252 336472
rect 284496 316006 284892 316034
rect 287072 316006 287468 316034
rect 288452 316006 288756 316034
rect 284496 294710 284524 316006
rect 284484 294704 284536 294710
rect 284484 294646 284536 294652
rect 287072 139398 287100 316006
rect 287060 139392 287112 139398
rect 287060 139334 287112 139340
rect 287060 54528 287112 54534
rect 287060 54470 287112 54476
rect 287072 16574 287100 54470
rect 288452 20670 288480 316006
rect 288440 20664 288492 20670
rect 288440 20606 288492 20612
rect 284404 16546 284984 16574
rect 287072 16546 287376 16574
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286600 5092 286652 5098
rect 286600 5034 286652 5040
rect 286612 480 286640 5034
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 291212 6914 291240 336466
rect 291304 7818 291332 338014
rect 292580 323604 292632 323610
rect 292580 323546 292632 323552
rect 291292 7812 291344 7818
rect 291292 7754 291344 7760
rect 291212 6886 291424 6914
rect 288992 4072 289044 4078
rect 288992 4014 289044 4020
rect 289004 480 289032 4014
rect 290188 4004 290240 4010
rect 290188 3946 290240 3952
rect 290200 480 290228 3946
rect 291396 480 291424 6886
rect 292592 480 292620 323546
rect 293236 316034 293264 338014
rect 294524 316034 294552 338014
rect 295812 316034 295840 338014
rect 296720 336456 296772 336462
rect 296720 336398 296772 336404
rect 292684 316006 293264 316034
rect 293972 316006 294552 316034
rect 295352 316006 295840 316034
rect 292684 280838 292712 316006
rect 292672 280832 292724 280838
rect 292672 280774 292724 280780
rect 293972 262886 294000 316006
rect 294052 263016 294104 263022
rect 294052 262958 294104 262964
rect 293960 262880 294012 262886
rect 293960 262822 294012 262828
rect 294064 16574 294092 262958
rect 295352 91798 295380 316006
rect 295340 91792 295392 91798
rect 295340 91734 295392 91740
rect 294064 16546 294920 16574
rect 293684 5976 293736 5982
rect 293684 5918 293736 5924
rect 293696 480 293724 5918
rect 294892 480 294920 16546
rect 296076 6112 296128 6118
rect 296076 6054 296128 6060
rect 296088 480 296116 6054
rect 296732 3482 296760 336398
rect 297100 316034 297128 338014
rect 298100 334892 298152 334898
rect 298100 334834 298152 334840
rect 296824 316006 297128 316034
rect 296824 6390 296852 316006
rect 296812 6384 296864 6390
rect 296812 6326 296864 6332
rect 296732 3454 297312 3482
rect 297284 480 297312 3454
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 334834
rect 298388 316034 298416 338014
rect 299676 316034 299704 338014
rect 300964 316034 300992 338014
rect 302238 336560 302294 336569
rect 302238 336495 302294 336504
rect 298204 316006 298416 316034
rect 299492 316006 299704 316034
rect 300872 316006 300992 316034
rect 298204 43450 298232 316006
rect 298192 43444 298244 43450
rect 298192 43386 298244 43392
rect 299492 6662 299520 316006
rect 300872 152522 300900 316006
rect 300860 152516 300912 152522
rect 300860 152458 300912 152464
rect 300768 9240 300820 9246
rect 300768 9182 300820 9188
rect 299480 6656 299532 6662
rect 299480 6598 299532 6604
rect 299664 3936 299716 3942
rect 299664 3878 299716 3884
rect 299676 480 299704 3878
rect 300780 480 300808 9182
rect 301964 8016 302016 8022
rect 301964 7958 302016 7964
rect 301976 480 302004 7958
rect 302252 3482 302280 336495
rect 302344 6390 302372 338014
rect 303620 331968 303672 331974
rect 303620 331910 303672 331916
rect 303632 16574 303660 331910
rect 303632 16546 303936 16574
rect 302332 6384 302384 6390
rect 302332 6326 302384 6332
rect 302252 3454 303200 3482
rect 303172 480 303200 3454
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305012 7886 305040 338014
rect 306392 246362 306420 338014
rect 307818 337770 307846 338028
rect 308692 338014 309120 338042
rect 309980 338014 310408 338042
rect 312004 338014 312340 338042
rect 313292 338014 313628 338042
rect 314672 338014 314916 338042
rect 316144 338014 316204 338042
rect 317432 338014 317492 338042
rect 318352 338014 318780 338042
rect 320928 338014 321356 338042
rect 322216 338014 322644 338042
rect 323596 338014 323932 338042
rect 324884 338014 325220 338042
rect 326080 338014 326508 338042
rect 327368 338014 327796 338042
rect 328656 338014 329084 338042
rect 329852 338014 330372 338042
rect 331876 338014 332304 338042
rect 333164 338014 333592 338042
rect 334452 338014 334880 338042
rect 335740 338014 336168 338042
rect 337028 338014 337456 338042
rect 338316 338014 338744 338042
rect 339604 338014 340032 338042
rect 341076 338014 341320 338042
rect 342608 338014 342944 338042
rect 307818 337742 307892 337770
rect 307760 331968 307812 331974
rect 307760 331910 307812 331916
rect 306380 246356 306432 246362
rect 306380 246298 306432 246304
rect 305000 7880 305052 7886
rect 305000 7822 305052 7828
rect 305552 7880 305604 7886
rect 305552 7822 305604 7828
rect 305564 480 305592 7822
rect 306748 6860 306800 6866
rect 306748 6802 306800 6808
rect 306760 480 306788 6802
rect 307772 2922 307800 331910
rect 307864 14482 307892 337742
rect 308692 316034 308720 338014
rect 309980 316034 310008 338014
rect 312004 333130 312032 338014
rect 311992 333124 312044 333130
rect 311992 333066 312044 333072
rect 311900 330608 311952 330614
rect 311900 330550 311952 330556
rect 310520 319592 310572 319598
rect 310520 319534 310572 319540
rect 307956 316006 308720 316034
rect 309152 316006 310008 316034
rect 307956 21418 307984 316006
rect 309152 296002 309180 316006
rect 309140 295996 309192 296002
rect 309140 295938 309192 295944
rect 307944 21412 307996 21418
rect 307944 21354 307996 21360
rect 310532 16574 310560 319534
rect 311912 16574 311940 330550
rect 313292 272542 313320 338014
rect 313280 272536 313332 272542
rect 313280 272478 313332 272484
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 307852 14476 307904 14482
rect 307852 14418 307904 14424
rect 310242 6624 310298 6633
rect 310242 6559 310298 6568
rect 307944 5160 307996 5166
rect 307944 5102 307996 5108
rect 307760 2916 307812 2922
rect 307760 2858 307812 2864
rect 307956 480 307984 5102
rect 309048 2916 309100 2922
rect 309048 2858 309100 2864
rect 309060 480 309088 2858
rect 310256 480 310284 6559
rect 311452 480 311480 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 314672 13122 314700 338014
rect 316038 336696 316094 336705
rect 316038 336631 316094 336640
rect 316052 16574 316080 336631
rect 316144 282198 316172 338014
rect 316132 282192 316184 282198
rect 316132 282134 316184 282140
rect 316052 16546 316264 16574
rect 314660 13116 314712 13122
rect 314660 13058 314712 13064
rect 313832 6792 313884 6798
rect 313832 6734 313884 6740
rect 313844 480 313872 6734
rect 315028 3596 315080 3602
rect 315028 3538 315080 3544
rect 315040 480 315068 3538
rect 316236 480 316264 16546
rect 317328 4956 317380 4962
rect 317328 4898 317380 4904
rect 317340 480 317368 4898
rect 317432 3534 317460 338014
rect 317512 330676 317564 330682
rect 317512 330618 317564 330624
rect 317524 16574 317552 330618
rect 318352 316034 318380 338014
rect 318798 337512 318854 337521
rect 318798 337447 318854 337456
rect 317616 316006 318380 316034
rect 317616 306338 317644 316006
rect 317604 306332 317656 306338
rect 317604 306274 317656 306280
rect 318812 16574 318840 337447
rect 320180 335708 320232 335714
rect 320180 335650 320232 335656
rect 320192 16574 320220 335650
rect 320928 316034 320956 338014
rect 322216 316034 322244 338014
rect 323596 336190 323624 338014
rect 323584 336184 323636 336190
rect 323584 336126 323636 336132
rect 324884 333946 324912 338014
rect 324872 333940 324924 333946
rect 324872 333882 324924 333888
rect 326080 316034 326108 338014
rect 327368 316034 327396 338014
rect 328656 316034 328684 338014
rect 329852 325650 329880 338014
rect 329840 325644 329892 325650
rect 329840 325586 329892 325592
rect 331876 316034 331904 338014
rect 333164 316034 333192 338014
rect 333980 337544 334032 337550
rect 333980 337486 334032 337492
rect 320284 316006 320956 316034
rect 321572 316006 322244 316034
rect 325712 316006 326108 316034
rect 327092 316006 327396 316034
rect 328472 316006 328684 316034
rect 331232 316006 331904 316034
rect 332612 316006 333192 316034
rect 320284 291854 320312 316006
rect 320272 291848 320324 291854
rect 320272 291790 320324 291796
rect 321572 47666 321600 316006
rect 324320 305720 324372 305726
rect 324320 305662 324372 305668
rect 322940 296064 322992 296070
rect 322940 296006 322992 296012
rect 321560 47660 321612 47666
rect 321560 47602 321612 47608
rect 317524 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 317420 3528 317472 3534
rect 317420 3470 317472 3476
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322112 6384 322164 6390
rect 322112 6326 322164 6332
rect 322124 480 322152 6326
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 296006
rect 324332 3534 324360 305662
rect 325712 22778 325740 316006
rect 325700 22772 325752 22778
rect 325700 22714 325752 22720
rect 326344 14476 326396 14482
rect 326344 14418 326396 14424
rect 324412 6588 324464 6594
rect 324412 6530 324464 6536
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 324424 480 324452 6530
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 14418
rect 327092 10334 327120 316006
rect 328472 257378 328500 316006
rect 329840 309800 329892 309806
rect 329840 309742 329892 309748
rect 328460 257372 328512 257378
rect 328460 257314 328512 257320
rect 329852 16574 329880 309742
rect 329852 16546 330432 16574
rect 327080 10328 327132 10334
rect 327080 10270 327132 10276
rect 327998 3904 328054 3913
rect 327998 3839 328054 3848
rect 328012 480 328040 3839
rect 329194 3224 329250 3233
rect 329194 3159 329250 3168
rect 329208 480 329236 3159
rect 330404 480 330432 16546
rect 331232 10334 331260 316006
rect 331312 123480 331364 123486
rect 331312 123422 331364 123428
rect 331220 10328 331272 10334
rect 331220 10270 331272 10276
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331324 354 331352 123422
rect 332612 5030 332640 316006
rect 332692 31068 332744 31074
rect 332692 31010 332744 31016
rect 332600 5024 332652 5030
rect 332600 4966 332652 4972
rect 332600 3868 332652 3874
rect 332600 3810 332652 3816
rect 332612 1986 332640 3810
rect 332704 3534 332732 31010
rect 333992 16574 334020 337486
rect 334452 316034 334480 338014
rect 335740 316034 335768 338014
rect 337028 316034 337056 338014
rect 338316 316034 338344 338014
rect 339604 316034 339632 338014
rect 340880 334892 340932 334898
rect 340880 334834 340932 334840
rect 334084 316006 334480 316034
rect 335372 316006 335768 316034
rect 336752 316006 337056 316034
rect 338132 316006 338344 316034
rect 339512 316006 339632 316034
rect 334084 46238 334112 316006
rect 334072 46232 334124 46238
rect 334072 46174 334124 46180
rect 333992 16546 334664 16574
rect 332692 3528 332744 3534
rect 332692 3470 332744 3476
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 332612 1958 332732 1986
rect 332704 480 332732 1958
rect 333900 480 333928 3470
rect 331558 354 331670 480
rect 331324 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 335372 6526 335400 316006
rect 335452 291916 335504 291922
rect 335452 291858 335504 291864
rect 335464 16574 335492 291858
rect 336752 25634 336780 316006
rect 338132 45558 338160 316006
rect 338120 45552 338172 45558
rect 338120 45494 338172 45500
rect 336740 25628 336792 25634
rect 336740 25570 336792 25576
rect 335464 16546 336320 16574
rect 335360 6520 335412 6526
rect 335360 6462 335412 6468
rect 336292 480 336320 16546
rect 339512 6730 339540 316006
rect 339500 6724 339552 6730
rect 339500 6666 339552 6672
rect 339868 5228 339920 5234
rect 339868 5170 339920 5176
rect 338672 4956 338724 4962
rect 338672 4898 338724 4904
rect 337474 4040 337530 4049
rect 337474 3975 337530 3984
rect 337488 480 337516 3975
rect 338684 480 338712 4898
rect 339880 480 339908 5170
rect 340892 3534 340920 334834
rect 340972 322312 341024 322318
rect 340972 322254 341024 322260
rect 340880 3528 340932 3534
rect 340880 3470 340932 3476
rect 340984 480 341012 322254
rect 341076 284986 341104 338014
rect 342916 336666 342944 338014
rect 343652 338014 343896 338042
rect 345124 338014 345184 338042
rect 346472 338014 346624 338042
rect 342904 336660 342956 336666
rect 342904 336602 342956 336608
rect 342260 336184 342312 336190
rect 342260 336126 342312 336132
rect 341064 284980 341116 284986
rect 341064 284922 341116 284928
rect 342272 16574 342300 336126
rect 343652 90370 343680 338014
rect 345020 309868 345072 309874
rect 345020 309810 345072 309816
rect 343640 90364 343692 90370
rect 343640 90306 343692 90312
rect 343640 25560 343692 25566
rect 343640 25502 343692 25508
rect 343652 16574 343680 25502
rect 345032 16574 345060 309810
rect 345124 303074 345152 338014
rect 346400 330472 346452 330478
rect 346400 330414 346452 330420
rect 345112 303068 345164 303074
rect 345112 303010 345164 303016
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 342180 480 342208 3470
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346412 7954 346440 330414
rect 346492 323672 346544 323678
rect 346492 323614 346544 323620
rect 346504 16574 346532 323614
rect 346596 303006 346624 338014
rect 347424 338014 347760 338042
rect 348620 338014 349048 338042
rect 350552 338014 350980 338042
rect 351932 338014 352268 338042
rect 353404 338014 353556 338042
rect 354692 338014 354844 338042
rect 356072 338014 356132 338042
rect 356992 338014 357420 338042
rect 358280 338014 358708 338042
rect 359568 338014 359996 338042
rect 360764 338014 361284 338042
rect 362144 338014 362572 338042
rect 363432 338014 363860 338042
rect 364720 338014 365148 338042
rect 366100 338014 366436 338042
rect 367296 338014 367724 338042
rect 368584 338014 369012 338042
rect 370516 338014 370944 338042
rect 371804 338014 372232 338042
rect 373092 338014 373520 338042
rect 374380 338014 374808 338042
rect 375668 338014 376096 338042
rect 376956 338014 377384 338042
rect 378336 338014 378672 338042
rect 347424 330478 347452 338014
rect 347780 333124 347832 333130
rect 347780 333066 347832 333072
rect 347412 330472 347464 330478
rect 347412 330414 347464 330420
rect 346584 303000 346636 303006
rect 346584 302942 346636 302948
rect 346504 16546 346992 16574
rect 346400 7948 346452 7954
rect 346400 7890 346452 7896
rect 346964 480 346992 16546
rect 347792 3482 347820 333066
rect 348620 316034 348648 338014
rect 349160 330676 349212 330682
rect 349160 330618 349212 330624
rect 347884 316006 348648 316034
rect 347884 5030 347912 316006
rect 349172 16574 349200 330618
rect 349172 16546 349292 16574
rect 347872 5024 347924 5030
rect 347872 4966 347924 4972
rect 347792 3454 348096 3482
rect 348068 480 348096 3454
rect 349264 480 349292 16546
rect 350552 5234 350580 338014
rect 350540 5228 350592 5234
rect 350540 5170 350592 5176
rect 351642 4040 351698 4049
rect 351642 3975 351698 3984
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 350460 480 350488 3470
rect 351656 480 351684 3975
rect 351932 3670 351960 338014
rect 352012 333056 352064 333062
rect 352012 332998 352064 333004
rect 352024 16574 352052 332998
rect 353300 325168 353352 325174
rect 353300 325110 353352 325116
rect 353312 16574 353340 325110
rect 353404 28286 353432 338014
rect 353392 28280 353444 28286
rect 353392 28222 353444 28228
rect 352024 16546 352880 16574
rect 353312 16546 353616 16574
rect 351920 3664 351972 3670
rect 351920 3606 351972 3612
rect 352852 480 352880 16546
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 354692 6594 354720 338014
rect 356072 333538 356100 338014
rect 356060 333532 356112 333538
rect 356060 333474 356112 333480
rect 356992 316034 357020 338014
rect 357440 336524 357492 336530
rect 357440 336466 357492 336472
rect 356072 316006 357020 316034
rect 354680 6588 354732 6594
rect 354680 6530 354732 6536
rect 356072 5166 356100 316006
rect 356334 6488 356390 6497
rect 356334 6423 356390 6432
rect 356060 5160 356112 5166
rect 356060 5102 356112 5108
rect 355232 3664 355284 3670
rect 355232 3606 355284 3612
rect 355244 480 355272 3606
rect 356348 480 356376 6423
rect 357452 3398 357480 336466
rect 358280 316034 358308 338014
rect 358818 337512 358874 337521
rect 358818 337447 358874 337456
rect 357544 316006 358308 316034
rect 357544 13122 357572 316006
rect 357532 13116 357584 13122
rect 357532 13058 357584 13064
rect 357532 6520 357584 6526
rect 357532 6462 357584 6468
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 6462
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 358832 626 358860 337447
rect 359568 316034 359596 338014
rect 360764 316034 360792 338014
rect 360936 335640 360988 335646
rect 360936 335582 360988 335588
rect 360948 316034 360976 335582
rect 362144 316034 362172 338014
rect 363432 316034 363460 338014
rect 364340 334960 364392 334966
rect 364340 334902 364392 334908
rect 358924 316006 359596 316034
rect 360212 316006 360792 316034
rect 360856 316006 360976 316034
rect 361592 316006 362172 316034
rect 363064 316006 363460 316034
rect 358924 5098 358952 316006
rect 360212 247722 360240 316006
rect 360200 247716 360252 247722
rect 360200 247658 360252 247664
rect 360856 65550 360884 316006
rect 361592 284986 361620 316006
rect 361580 284980 361632 284986
rect 361580 284922 361632 284928
rect 360844 65544 360896 65550
rect 360844 65486 360896 65492
rect 362316 9172 362368 9178
rect 362316 9114 362368 9120
rect 361120 6384 361172 6390
rect 361120 6326 361172 6332
rect 358912 5092 358964 5098
rect 358912 5034 358964 5040
rect 358832 598 359504 626
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 598
rect 361132 480 361160 6326
rect 362328 480 362356 9114
rect 363064 3505 363092 316006
rect 363512 6452 363564 6458
rect 363512 6394 363564 6400
rect 363050 3496 363106 3505
rect 363050 3431 363106 3440
rect 363524 480 363552 6394
rect 364352 3482 364380 334902
rect 364720 316034 364748 338014
rect 366100 335646 366128 338014
rect 367100 336592 367152 336598
rect 367100 336534 367152 336540
rect 366088 335640 366140 335646
rect 366088 335582 366140 335588
rect 364444 316006 364748 316034
rect 364444 3641 364472 316006
rect 365720 86284 365772 86290
rect 365720 86226 365772 86232
rect 364430 3632 364486 3641
rect 364430 3567 364486 3576
rect 364352 3454 364656 3482
rect 364628 480 364656 3454
rect 365732 3398 365760 86226
rect 367112 6914 367140 336534
rect 367296 316034 367324 338014
rect 367742 337376 367798 337385
rect 367742 337311 367798 337320
rect 367204 316006 367324 316034
rect 367204 17270 367232 316006
rect 367192 17264 367244 17270
rect 367192 17206 367244 17212
rect 367756 16574 367784 337311
rect 368584 316034 368612 338014
rect 370516 316034 370544 338014
rect 371804 316034 371832 338014
rect 373092 316034 373120 338014
rect 374000 333532 374052 333538
rect 374000 333474 374052 333480
rect 368492 316006 368612 316034
rect 369964 316006 370544 316034
rect 371252 316006 371832 316034
rect 372632 316006 373120 316034
rect 368492 25566 368520 316006
rect 369860 308508 369912 308514
rect 369860 308450 369912 308456
rect 368572 57248 368624 57254
rect 368572 57190 368624 57196
rect 368480 25560 368532 25566
rect 368480 25502 368532 25508
rect 368584 16574 368612 57190
rect 369872 16574 369900 308450
rect 369964 268462 369992 316006
rect 369952 268456 370004 268462
rect 369952 268398 370004 268404
rect 367756 16546 367876 16574
rect 368584 16546 369440 16574
rect 369872 16546 370176 16574
rect 367112 6886 367784 6914
rect 365810 6488 365866 6497
rect 365810 6423 365866 6432
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 480 365852 6423
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 6886
rect 367848 3874 367876 16546
rect 367836 3868 367888 3874
rect 367836 3810 367888 3816
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 371252 15910 371280 316006
rect 371240 15904 371292 15910
rect 371240 15846 371292 15852
rect 372632 4826 372660 316006
rect 372712 32428 372764 32434
rect 372712 32370 372764 32376
rect 372724 16574 372752 32370
rect 374012 16574 374040 333474
rect 374380 316034 374408 338014
rect 375380 334824 375432 334830
rect 375380 334766 375432 334772
rect 374104 316006 374408 316034
rect 374104 305726 374132 316006
rect 374092 305720 374144 305726
rect 374092 305662 374144 305668
rect 375392 16574 375420 334766
rect 375668 316034 375696 338014
rect 376760 337612 376812 337618
rect 376760 337554 376812 337560
rect 375484 316006 375696 316034
rect 375484 268394 375512 316006
rect 375472 268388 375524 268394
rect 375472 268330 375524 268336
rect 376772 16574 376800 337554
rect 376956 316034 376984 338014
rect 378336 336734 378364 338014
rect 378324 336728 378376 336734
rect 378324 336670 378376 336676
rect 378784 336728 378836 336734
rect 378784 336670 378836 336676
rect 376864 316006 376984 316034
rect 376864 206990 376892 316006
rect 378140 282192 378192 282198
rect 378140 282134 378192 282140
rect 376852 206984 376904 206990
rect 376852 206926 376904 206932
rect 378152 16574 378180 282134
rect 378796 69698 378824 336670
rect 378784 69692 378836 69698
rect 378784 69634 378836 69640
rect 372724 16546 372936 16574
rect 374012 16546 374132 16574
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 372620 4820 372672 4826
rect 372620 4762 372672 4768
rect 371700 3800 371752 3806
rect 371700 3742 371752 3748
rect 371712 480 371740 3742
rect 372908 480 372936 16546
rect 374104 480 374132 16546
rect 375288 6452 375340 6458
rect 375288 6394 375340 6400
rect 375300 480 375328 6394
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 370566 -960 370678 326
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 338127
rect 379624 338014 379960 338042
rect 380912 338014 381248 338042
rect 382476 338014 382536 338042
rect 383764 338014 383824 338042
rect 385052 338014 385112 338042
rect 385972 338014 386400 338042
rect 387260 338014 387688 338042
rect 389284 338014 389620 338042
rect 390572 338014 390908 338042
rect 391952 338014 392196 338042
rect 393332 338014 393484 338042
rect 394772 338014 394924 338042
rect 379624 24138 379652 338014
rect 380912 336734 380940 338014
rect 380900 336728 380952 336734
rect 380900 336670 380952 336676
rect 381544 335980 381596 335986
rect 381544 335922 381596 335928
rect 380992 335640 381044 335646
rect 380992 335582 381044 335588
rect 379612 24132 379664 24138
rect 379612 24074 379664 24080
rect 381004 16574 381032 335582
rect 381004 16546 381216 16574
rect 381188 480 381216 16546
rect 381556 3369 381584 335922
rect 382280 330540 382332 330546
rect 382280 330482 382332 330488
rect 381542 3360 381598 3369
rect 381542 3295 381598 3304
rect 382292 3210 382320 330482
rect 382370 316976 382426 316985
rect 382370 316911 382426 316920
rect 382384 3398 382412 316911
rect 382476 235278 382504 338014
rect 383660 326528 383712 326534
rect 383660 326470 383712 326476
rect 382464 235272 382516 235278
rect 382464 235214 382516 235220
rect 383672 16574 383700 326470
rect 383764 64190 383792 338014
rect 385052 150414 385080 338014
rect 385972 316034 386000 338014
rect 387260 316742 387288 338014
rect 387800 337680 387852 337686
rect 387800 337622 387852 337628
rect 387248 316736 387300 316742
rect 387248 316678 387300 316684
rect 385144 316006 386000 316034
rect 385144 269822 385172 316006
rect 385132 269816 385184 269822
rect 385132 269758 385184 269764
rect 386420 233980 386472 233986
rect 386420 233922 386472 233928
rect 385040 150408 385092 150414
rect 385040 150350 385092 150356
rect 383752 64184 383804 64190
rect 383752 64126 383804 64132
rect 386432 16574 386460 233922
rect 383672 16546 384344 16574
rect 386432 16546 386736 16574
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382292 3182 382412 3210
rect 382384 480 382412 3182
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385960 6588 386012 6594
rect 385960 6530 386012 6536
rect 385972 480 386000 6530
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 337622
rect 389284 335986 389312 338014
rect 389272 335980 389324 335986
rect 389272 335922 389324 335928
rect 390572 333198 390600 338014
rect 390560 333192 390612 333198
rect 390560 333134 390612 333140
rect 390558 326360 390614 326369
rect 390558 326295 390614 326304
rect 389180 305720 389232 305726
rect 389180 305662 389232 305668
rect 389192 16574 389220 305662
rect 390572 16574 390600 326295
rect 389192 16546 389496 16574
rect 390572 16546 390692 16574
rect 389468 480 389496 16546
rect 390664 480 390692 16546
rect 391952 6458 391980 338014
rect 392032 17264 392084 17270
rect 392032 17206 392084 17212
rect 392044 16574 392072 17206
rect 392044 16546 392624 16574
rect 391940 6452 391992 6458
rect 391940 6394 391992 6400
rect 391846 3496 391902 3505
rect 391846 3431 391902 3440
rect 391860 480 391888 3431
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 393332 6186 393360 338014
rect 394700 337748 394752 337754
rect 394700 337690 394752 337696
rect 393412 319524 393464 319530
rect 393412 319466 393464 319472
rect 393424 16574 393452 319466
rect 394712 16574 394740 337690
rect 394792 326800 394844 326806
rect 394792 326742 394844 326748
rect 394804 24138 394832 326742
rect 394896 303006 394924 338014
rect 395724 338014 396060 338042
rect 397288 338014 397348 338042
rect 398636 338014 398788 338042
rect 395724 326806 395752 338014
rect 397288 333810 397316 338014
rect 398760 333946 398788 338014
rect 398944 335354 398972 338127
rect 398852 335326 398972 335354
rect 399496 338014 399924 338042
rect 400784 338014 401212 338042
rect 402164 338014 402500 338042
rect 405076 338014 405412 338042
rect 398748 333940 398800 333946
rect 398748 333882 398800 333888
rect 397276 333804 397328 333810
rect 397276 333746 397328 333752
rect 395712 326800 395764 326806
rect 395712 326742 395764 326748
rect 394884 303000 394936 303006
rect 394884 302942 394936 302948
rect 396080 280832 396132 280838
rect 396080 280774 396132 280780
rect 394792 24132 394844 24138
rect 394792 24074 394844 24080
rect 393424 16546 394280 16574
rect 394712 16546 395384 16574
rect 393320 6180 393372 6186
rect 393320 6122 393372 6128
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 280774
rect 397460 60036 397512 60042
rect 397460 59978 397512 59984
rect 397472 16574 397500 59978
rect 398852 16574 398880 335326
rect 399496 316034 399524 338014
rect 400220 329112 400272 329118
rect 400220 329054 400272 329060
rect 398944 316006 399524 316034
rect 398944 39370 398972 316006
rect 398932 39364 398984 39370
rect 398932 39306 398984 39312
rect 400232 16574 400260 329054
rect 400784 316034 400812 338014
rect 402164 336734 402192 338014
rect 400864 336728 400916 336734
rect 400864 336670 400916 336676
rect 402152 336728 402204 336734
rect 402152 336670 402204 336676
rect 400324 316006 400812 316034
rect 400324 305726 400352 316006
rect 400312 305720 400364 305726
rect 400312 305662 400364 305668
rect 400876 51746 400904 336670
rect 405384 335986 405412 338014
rect 405936 338014 406364 338042
rect 407224 338014 407652 338042
rect 409156 338014 409584 338042
rect 410444 338014 410872 338042
rect 413112 338014 413448 338042
rect 414308 338014 414736 338042
rect 415596 338014 416024 338042
rect 416976 338014 417312 338042
rect 418264 338014 418600 338042
rect 419888 338014 420224 338042
rect 405740 337816 405792 337822
rect 405740 337758 405792 337764
rect 405372 335980 405424 335986
rect 405372 335922 405424 335928
rect 405004 335844 405056 335850
rect 405004 335786 405056 335792
rect 402980 303068 403032 303074
rect 402980 303010 403032 303016
rect 400864 51740 400916 51746
rect 400864 51682 400916 51688
rect 402992 16574 403020 303010
rect 405016 55894 405044 335786
rect 405004 55888 405056 55894
rect 405004 55830 405056 55836
rect 405752 16574 405780 337758
rect 405936 316034 405964 338014
rect 407120 335912 407172 335918
rect 407120 335854 407172 335860
rect 405844 316006 405964 316034
rect 405844 233918 405872 316006
rect 405832 233912 405884 233918
rect 405832 233854 405884 233860
rect 397472 16546 397776 16574
rect 398852 16546 398972 16574
rect 400232 16546 400904 16574
rect 402992 16546 403664 16574
rect 405752 16546 406056 16574
rect 397748 480 397776 16546
rect 398944 480 398972 16546
rect 400128 9104 400180 9110
rect 400128 9046 400180 9052
rect 400140 480 400168 9046
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402520 5024 402572 5030
rect 402520 4966 402572 4972
rect 402532 480 402560 4966
rect 403636 480 403664 16546
rect 404820 3800 404872 3806
rect 404820 3742 404872 3748
rect 404832 480 404860 3742
rect 406028 480 406056 16546
rect 407132 3398 407160 335854
rect 407224 16574 407252 338014
rect 409156 316034 409184 338014
rect 409880 337952 409932 337958
rect 409880 337894 409932 337900
rect 408512 316006 409184 316034
rect 407224 16546 407344 16574
rect 407212 6248 407264 6254
rect 407212 6190 407264 6196
rect 407120 3392 407172 3398
rect 407120 3334 407172 3340
rect 407224 480 407252 6190
rect 407316 4894 407344 16546
rect 408512 6526 408540 316006
rect 408592 300144 408644 300150
rect 408592 300086 408644 300092
rect 408604 16574 408632 300086
rect 408604 16546 409184 16574
rect 408500 6520 408552 6526
rect 408500 6462 408552 6468
rect 407304 4888 407356 4894
rect 407304 4830 407356 4836
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 409892 3482 409920 337894
rect 410444 316034 410472 338014
rect 413112 336122 413140 338014
rect 413100 336116 413152 336122
rect 413100 336058 413152 336064
rect 414308 316034 414336 338014
rect 415400 334824 415452 334830
rect 415400 334766 415452 334772
rect 409984 316006 410472 316034
rect 414032 316006 414336 316034
rect 409984 4962 410012 316006
rect 411260 256012 411312 256018
rect 411260 255954 411312 255960
rect 411272 16574 411300 255954
rect 411272 16546 411944 16574
rect 409972 4956 410024 4962
rect 409972 4898 410024 4904
rect 409892 3454 410840 3482
rect 410812 480 410840 3454
rect 411916 480 411944 16546
rect 414032 4894 414060 316006
rect 415412 6914 415440 334766
rect 415596 316034 415624 338014
rect 416976 336054 417004 338014
rect 416964 336048 417016 336054
rect 416964 335990 417016 335996
rect 418160 333804 418212 333810
rect 418160 333746 418212 333752
rect 415504 316006 415624 316034
rect 415504 7750 415532 316006
rect 416780 80708 416832 80714
rect 416780 80650 416832 80656
rect 416792 16574 416820 80650
rect 418172 16574 418200 333746
rect 418264 17270 418292 338014
rect 419540 337884 419592 337890
rect 419540 337826 419592 337832
rect 418252 17264 418304 17270
rect 418252 17206 418304 17212
rect 419552 16574 419580 337826
rect 420196 336054 420224 338014
rect 421024 338014 421176 338042
rect 422312 338014 422464 338042
rect 423692 338014 423752 338042
rect 424980 338014 425040 338042
rect 425992 338014 426328 338042
rect 427924 338014 428260 338042
rect 429304 338014 429548 338042
rect 430684 338014 430836 338042
rect 431972 338014 432124 338042
rect 433352 338014 433412 338042
rect 434272 338014 434700 338042
rect 435560 338014 435988 338042
rect 436664 338014 437276 338042
rect 438136 338014 438564 338042
rect 439424 338014 439852 338042
rect 441140 338014 441384 338042
rect 420184 336048 420236 336054
rect 420184 335990 420236 335996
rect 420920 322244 420972 322250
rect 420920 322186 420972 322192
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 415492 7744 415544 7750
rect 415492 7686 415544 7692
rect 415412 6886 415532 6914
rect 414020 4888 414072 4894
rect 414020 4830 414072 4836
rect 413100 4820 413152 4826
rect 413100 4762 413152 4768
rect 413112 480 413140 4762
rect 414296 4004 414348 4010
rect 414296 3946 414348 3952
rect 414308 480 414336 3946
rect 415504 480 415532 6886
rect 416688 3936 416740 3942
rect 416688 3878 416740 3884
rect 416700 480 416728 3878
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 322186
rect 421024 18630 421052 338014
rect 421012 18624 421064 18630
rect 421012 18566 421064 18572
rect 422312 4214 422340 338014
rect 423692 336734 423720 338014
rect 422944 336728 422996 336734
rect 422944 336670 422996 336676
rect 423680 336728 423732 336734
rect 423680 336670 423732 336676
rect 422392 254584 422444 254590
rect 422392 254526 422444 254532
rect 422404 16574 422432 254526
rect 422956 250510 422984 336670
rect 424980 336122 425008 338014
rect 424968 336116 425020 336122
rect 424968 336058 425020 336064
rect 425992 335850 426020 338014
rect 427924 336734 427952 338014
rect 428004 337340 428056 337346
rect 428004 337282 428056 337288
rect 427084 336728 427136 336734
rect 427084 336670 427136 336676
rect 427912 336728 427964 336734
rect 427912 336670 427964 336676
rect 425980 335844 426032 335850
rect 425980 335786 426032 335792
rect 427096 263022 427124 336670
rect 428016 316034 428044 337282
rect 429200 333192 429252 333198
rect 429200 333134 429252 333140
rect 427924 316006 428044 316034
rect 427084 263016 427136 263022
rect 427084 262958 427136 262964
rect 422944 250504 422996 250510
rect 422944 250446 422996 250452
rect 423680 173188 423732 173194
rect 423680 173130 423732 173136
rect 422404 16546 422616 16574
rect 422300 4208 422352 4214
rect 422300 4150 422352 4156
rect 422588 480 422616 16546
rect 423692 3398 423720 173130
rect 427924 16574 427952 316006
rect 427924 16546 428504 16574
rect 426164 8968 426216 8974
rect 426164 8910 426216 8916
rect 423772 4208 423824 4214
rect 423772 4150 423824 4156
rect 423680 3392 423732 3398
rect 423680 3334 423732 3340
rect 423784 480 423812 4150
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 426176 480 426204 8910
rect 427268 4072 427320 4078
rect 427268 4014 427320 4020
rect 427280 480 427308 4014
rect 428476 480 428504 16546
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429212 354 429240 333134
rect 429304 6390 429332 338014
rect 430580 337272 430632 337278
rect 430580 337214 430632 337220
rect 429292 6384 429344 6390
rect 429292 6326 429344 6332
rect 430592 3482 430620 337214
rect 430684 6322 430712 338014
rect 431972 164898 432000 338014
rect 433352 335918 433380 338014
rect 433340 335912 433392 335918
rect 433340 335854 433392 335860
rect 434272 316034 434300 338014
rect 434720 337204 434772 337210
rect 434720 337146 434772 337152
rect 433444 316006 434300 316034
rect 433444 305726 433472 316006
rect 433432 305720 433484 305726
rect 433432 305662 433484 305668
rect 431960 164892 432012 164898
rect 431960 164834 432012 164840
rect 434732 16574 434760 337146
rect 435560 316034 435588 338014
rect 436664 316034 436692 338014
rect 436744 336048 436796 336054
rect 436744 335990 436796 335996
rect 434824 316006 435588 316034
rect 436112 316006 436692 316034
rect 434824 54534 434852 316006
rect 436112 308514 436140 316006
rect 436100 308508 436152 308514
rect 436100 308450 436152 308456
rect 434812 54528 434864 54534
rect 434812 54470 434864 54476
rect 434732 16546 435128 16574
rect 430672 6316 430724 6322
rect 430672 6258 430724 6264
rect 432052 4888 432104 4894
rect 432052 4830 432104 4836
rect 430592 3454 430896 3482
rect 430868 480 430896 3454
rect 432064 480 432092 4830
rect 434444 4140 434496 4146
rect 434444 4082 434496 4088
rect 433248 3120 433300 3126
rect 433248 3062 433300 3068
rect 433260 480 433288 3062
rect 434456 480 434484 4082
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 436756 5574 436784 335990
rect 438136 316034 438164 338014
rect 438860 334688 438912 334694
rect 438860 334630 438912 334636
rect 437492 316006 438164 316034
rect 437492 309874 437520 316006
rect 437480 309868 437532 309874
rect 437480 309810 437532 309816
rect 438872 16574 438900 334630
rect 439424 316034 439452 338014
rect 441356 336462 441384 338014
rect 442000 338014 442428 338042
rect 443288 338014 443716 338042
rect 444576 338014 445004 338042
rect 446292 338014 446628 338042
rect 441344 336456 441396 336462
rect 441344 336398 441396 336404
rect 440240 336048 440292 336054
rect 440240 335990 440292 335996
rect 438964 316006 439452 316034
rect 438964 289134 438992 316006
rect 438952 289128 439004 289134
rect 438952 289070 439004 289076
rect 440252 16574 440280 335990
rect 441618 334112 441674 334121
rect 441618 334047 441674 334056
rect 438872 16546 439176 16574
rect 440252 16546 440372 16574
rect 436744 5568 436796 5574
rect 436744 5510 436796 5516
rect 436742 3632 436798 3641
rect 436742 3567 436798 3576
rect 436756 480 436784 3567
rect 437938 3224 437994 3233
rect 437938 3159 437994 3168
rect 437952 480 437980 3159
rect 439148 480 439176 16546
rect 440344 480 440372 16546
rect 441632 6914 441660 334047
rect 442000 316034 442028 338014
rect 443288 316034 443316 338014
rect 444576 316034 444604 338014
rect 446600 336734 446628 338014
rect 446588 336728 446640 336734
rect 446588 336670 446640 336676
rect 441724 316006 442028 316034
rect 443012 316006 443316 316034
rect 444392 316006 444604 316034
rect 441724 7886 441752 316006
rect 441712 7880 441764 7886
rect 441712 7822 441764 7828
rect 443012 7614 443040 316006
rect 443000 7608 443052 7614
rect 443000 7550 443052 7556
rect 441632 6886 442672 6914
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 6886
rect 443828 5568 443880 5574
rect 443828 5510 443880 5516
rect 443840 480 443868 5510
rect 444392 4826 444420 316006
rect 445758 304192 445814 304201
rect 445758 304127 445814 304136
rect 444472 17264 444524 17270
rect 444472 17206 444524 17212
rect 444484 16574 444512 17206
rect 444484 16546 445064 16574
rect 444380 4820 444432 4826
rect 444380 4762 444432 4768
rect 445036 480 445064 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 304127
rect 447152 16574 447180 338166
rect 450358 338127 450414 338136
rect 447796 338014 448224 338042
rect 449084 338014 449512 338042
rect 447796 316034 447824 338014
rect 448520 337476 448572 337482
rect 448520 337418 448572 337424
rect 448532 335986 448560 337418
rect 448520 335980 448572 335986
rect 448520 335922 448572 335928
rect 449084 316034 449112 338014
rect 449898 337648 449954 337657
rect 449898 337583 449954 337592
rect 449164 336728 449216 336734
rect 449164 336670 449216 336676
rect 447244 316006 447824 316034
rect 448532 316006 449112 316034
rect 447244 215286 447272 316006
rect 448532 315314 448560 316006
rect 449176 315382 449204 336670
rect 449912 325038 449940 337583
rect 450372 335354 450400 338127
rect 450464 338014 450800 338042
rect 450464 336734 450492 338014
rect 451280 337136 451332 337142
rect 451280 337078 451332 337084
rect 450452 336728 450504 336734
rect 450452 336670 450504 336676
rect 450372 335326 450584 335354
rect 449900 325032 449952 325038
rect 449900 324974 449952 324980
rect 449164 315376 449216 315382
rect 449164 315318 449216 315324
rect 448520 315308 448572 315314
rect 448520 315250 448572 315256
rect 447782 293176 447838 293185
rect 447782 293111 447838 293120
rect 447232 215280 447284 215286
rect 447232 215222 447284 215228
rect 447152 16546 447456 16574
rect 446404 3596 446456 3602
rect 446404 3538 446456 3544
rect 446416 3330 446444 3538
rect 446404 3324 446456 3330
rect 446404 3266 446456 3272
rect 447428 480 447456 16546
rect 447796 3602 447824 293111
rect 450556 3738 450584 335326
rect 451292 16574 451320 337078
rect 451568 333062 451596 556990
rect 451660 555490 451688 559098
rect 451648 555484 451700 555490
rect 451648 555426 451700 555432
rect 451752 554062 451780 559846
rect 451740 554056 451792 554062
rect 451740 553998 451792 554004
rect 451646 513496 451702 513505
rect 451646 513431 451702 513440
rect 451660 333538 451688 513431
rect 451738 495136 451794 495145
rect 451738 495071 451794 495080
rect 451752 334830 451780 495071
rect 452672 491065 452700 670686
rect 453120 577516 453172 577522
rect 453120 577458 453172 577464
rect 453028 570716 453080 570722
rect 453028 570658 453080 570664
rect 452934 559872 452990 559881
rect 452934 559807 452990 559816
rect 452750 555112 452806 555121
rect 452750 555047 452806 555056
rect 452658 491056 452714 491065
rect 452658 490991 452714 491000
rect 451830 480176 451886 480185
rect 451830 480111 451886 480120
rect 451844 335714 451872 480111
rect 452106 474056 452162 474065
rect 452106 473991 452162 474000
rect 452014 457736 452070 457745
rect 452014 457671 452070 457680
rect 451924 355156 451976 355162
rect 451924 355098 451976 355104
rect 451832 335708 451884 335714
rect 451832 335650 451884 335656
rect 451740 334824 451792 334830
rect 451740 334766 451792 334772
rect 451648 333532 451700 333538
rect 451648 333474 451700 333480
rect 451556 333056 451608 333062
rect 451556 332998 451608 333004
rect 451292 16546 451688 16574
rect 450544 3732 450596 3738
rect 450544 3674 450596 3680
rect 447784 3596 447836 3602
rect 447784 3538 447836 3544
rect 448612 3596 448664 3602
rect 448612 3538 448664 3544
rect 448624 480 448652 3538
rect 449808 3256 449860 3262
rect 449808 3198 449860 3204
rect 449820 480 449848 3198
rect 450912 3188 450964 3194
rect 450912 3130 450964 3136
rect 450924 480 450952 3130
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 451936 3126 451964 355098
rect 452028 337550 452056 457671
rect 452016 337544 452068 337550
rect 452016 337486 452068 337492
rect 452120 334898 452148 473991
rect 452658 468616 452714 468625
rect 452658 468551 452660 468560
rect 452712 468551 452714 468560
rect 452660 468522 452712 468528
rect 452658 459096 452714 459105
rect 452658 459031 452714 459040
rect 452672 458454 452700 459031
rect 452660 458448 452712 458454
rect 452660 458390 452712 458396
rect 452764 430545 452792 555047
rect 452948 551342 452976 559807
rect 452936 551336 452988 551342
rect 452936 551278 452988 551284
rect 452842 531856 452898 531865
rect 452842 531791 452898 531800
rect 452750 430536 452806 430545
rect 452750 430471 452806 430480
rect 452752 425060 452804 425066
rect 452752 425002 452804 425008
rect 452764 423745 452792 425002
rect 452750 423736 452806 423745
rect 452750 423671 452806 423680
rect 452856 410009 452884 531791
rect 452936 523728 452988 523734
rect 452936 523670 452988 523676
rect 452842 410000 452898 410009
rect 452842 409935 452898 409944
rect 452658 409456 452714 409465
rect 452658 409391 452714 409400
rect 452672 408882 452700 409391
rect 452660 408876 452712 408882
rect 452660 408818 452712 408824
rect 452658 401296 452714 401305
rect 452658 401231 452714 401240
rect 452672 400246 452700 401231
rect 452660 400240 452712 400246
rect 452660 400182 452712 400188
rect 452198 391096 452254 391105
rect 452198 391031 452254 391040
rect 452212 337958 452240 391031
rect 452842 388376 452898 388385
rect 452842 388311 452898 388320
rect 452750 374776 452806 374785
rect 452750 374711 452806 374720
rect 452658 355056 452714 355065
rect 452658 354991 452714 355000
rect 452568 348832 452620 348838
rect 452568 348774 452620 348780
rect 452580 345014 452608 348774
rect 452304 344986 452608 345014
rect 452200 337952 452252 337958
rect 452200 337894 452252 337900
rect 452108 334892 452160 334898
rect 452108 334834 452160 334840
rect 452304 333130 452332 344986
rect 452384 342372 452436 342378
rect 452384 342314 452436 342320
rect 452292 333124 452344 333130
rect 452292 333066 452344 333072
rect 452396 3330 452424 342314
rect 452672 334762 452700 354991
rect 452660 334756 452712 334762
rect 452660 334698 452712 334704
rect 452764 87650 452792 374711
rect 452856 180130 452884 388311
rect 452948 355162 452976 523670
rect 453040 451625 453068 570658
rect 453132 514078 453160 577458
rect 453212 566500 453264 566506
rect 453212 566442 453264 566448
rect 453120 514072 453172 514078
rect 453120 514014 453172 514020
rect 453224 508065 453252 566442
rect 456984 562352 457036 562358
rect 456984 562294 457036 562300
rect 456892 559360 456944 559366
rect 456892 559302 456944 559308
rect 453304 558272 453356 558278
rect 453304 558214 453356 558220
rect 453210 508056 453266 508065
rect 453210 507991 453266 508000
rect 453210 482896 453266 482905
rect 453210 482831 453266 482840
rect 453224 482798 453252 482831
rect 453212 482792 453264 482798
rect 453212 482734 453264 482740
rect 453210 464536 453266 464545
rect 453210 464471 453266 464480
rect 453224 464234 453252 464471
rect 453212 464228 453264 464234
rect 453212 464170 453264 464176
rect 453026 451616 453082 451625
rect 453026 451551 453082 451560
rect 453026 447536 453082 447545
rect 453026 447471 453028 447480
rect 453080 447471 453082 447480
rect 453028 447442 453080 447448
rect 453026 427816 453082 427825
rect 453026 427751 453082 427760
rect 452936 355156 452988 355162
rect 452936 355098 452988 355104
rect 452934 344856 452990 344865
rect 452934 344791 452990 344800
rect 452948 343942 452976 344791
rect 452936 343936 452988 343942
rect 452936 343878 452988 343884
rect 453040 331906 453068 427751
rect 453210 416936 453266 416945
rect 453210 416871 453212 416880
rect 453264 416871 453266 416880
rect 453212 416842 453264 416848
rect 453210 382936 453266 382945
rect 453210 382871 453212 382880
rect 453264 382871 453266 382880
rect 453212 382842 453264 382848
rect 453118 380216 453174 380225
rect 453118 380151 453174 380160
rect 453028 331900 453080 331906
rect 453028 331842 453080 331848
rect 453132 308446 453160 380151
rect 453316 347750 453344 558214
rect 453580 557116 453632 557122
rect 453580 557058 453632 557064
rect 453394 550216 453450 550225
rect 453394 550151 453450 550160
rect 453408 549506 453436 550151
rect 453396 549500 453448 549506
rect 453396 549442 453448 549448
rect 453592 549250 453620 557058
rect 453672 556572 453724 556578
rect 453672 556514 453724 556520
rect 453408 549222 453620 549250
rect 453408 350402 453436 549222
rect 453684 547874 453712 556514
rect 454040 554804 454092 554810
rect 454040 554746 454092 554752
rect 453946 554296 454002 554305
rect 453946 554231 454002 554240
rect 453960 553450 453988 554231
rect 453948 553444 454000 553450
rect 453948 553386 454000 553392
rect 453500 547846 453712 547874
rect 453500 356046 453528 547846
rect 453946 547496 454002 547505
rect 453946 547431 454002 547440
rect 453960 546582 453988 547431
rect 453948 546576 454000 546582
rect 453948 546518 454000 546524
rect 453946 546136 454002 546145
rect 453946 546071 454002 546080
rect 453960 545154 453988 546071
rect 453948 545148 454000 545154
rect 453948 545090 454000 545096
rect 453578 544776 453634 544785
rect 453578 544711 453634 544720
rect 453592 544066 453620 544711
rect 453580 544060 453632 544066
rect 453580 544002 453632 544008
rect 453946 543416 454002 543425
rect 453946 543351 454002 543360
rect 453960 542434 453988 543351
rect 453948 542428 454000 542434
rect 453948 542370 454000 542376
rect 453762 542056 453818 542065
rect 453762 541991 453818 542000
rect 453776 541006 453804 541991
rect 453764 541000 453816 541006
rect 453764 540942 453816 540948
rect 453762 537976 453818 537985
rect 453762 537911 453818 537920
rect 453776 536858 453804 537911
rect 453764 536852 453816 536858
rect 453764 536794 453816 536800
rect 453946 535936 454002 535945
rect 453946 535871 454002 535880
rect 453960 535498 453988 535871
rect 453948 535492 454000 535498
rect 453948 535434 454000 535440
rect 453946 533216 454002 533225
rect 453946 533151 454002 533160
rect 453960 532778 453988 533151
rect 453948 532772 454000 532778
rect 453948 532714 454000 532720
rect 453578 530496 453634 530505
rect 453578 530431 453634 530440
rect 453592 523734 453620 530431
rect 453946 527776 454002 527785
rect 453946 527711 454002 527720
rect 453960 527202 453988 527711
rect 453948 527196 454000 527202
rect 453948 527138 454000 527144
rect 453670 525056 453726 525065
rect 453670 524991 453726 525000
rect 453684 524754 453712 524991
rect 453672 524748 453724 524754
rect 453672 524690 453724 524696
rect 453580 523728 453632 523734
rect 453580 523670 453632 523676
rect 453946 522336 454002 522345
rect 453946 522271 454002 522280
rect 453960 521694 453988 522271
rect 453948 521688 454000 521694
rect 453948 521630 454000 521636
rect 453946 520976 454002 520985
rect 453946 520911 453948 520920
rect 454000 520911 454002 520920
rect 453948 520882 454000 520888
rect 453946 519616 454002 519625
rect 453946 519551 454002 519560
rect 453960 518974 453988 519551
rect 453948 518968 454000 518974
rect 453948 518910 454000 518916
rect 453946 514856 454002 514865
rect 453946 514791 453948 514800
rect 454000 514791 454002 514800
rect 453948 514762 454000 514768
rect 453580 514072 453632 514078
rect 453580 514014 453632 514020
rect 453592 502625 453620 514014
rect 453764 513324 453816 513330
rect 453764 513266 453816 513272
rect 453776 512145 453804 513266
rect 453762 512136 453818 512145
rect 453762 512071 453818 512080
rect 453762 509416 453818 509425
rect 453762 509351 453818 509360
rect 453776 509318 453804 509351
rect 453764 509312 453816 509318
rect 453764 509254 453816 509260
rect 453946 503976 454002 503985
rect 453946 503911 454002 503920
rect 453960 503742 453988 503911
rect 453948 503736 454000 503742
rect 453948 503678 454000 503684
rect 453578 502616 453634 502625
rect 453578 502551 453634 502560
rect 453946 499896 454002 499905
rect 453946 499831 454002 499840
rect 453960 499594 453988 499831
rect 453948 499588 454000 499594
rect 453948 499530 454000 499536
rect 453946 498536 454002 498545
rect 453946 498471 453948 498480
rect 454000 498471 454002 498480
rect 453948 498442 454000 498448
rect 453948 492652 454000 492658
rect 453948 492594 454000 492600
rect 453960 492425 453988 492594
rect 453946 492416 454002 492425
rect 453946 492351 454002 492360
rect 453762 489696 453818 489705
rect 453762 489631 453818 489640
rect 453776 488578 453804 489631
rect 453764 488572 453816 488578
rect 453764 488514 453816 488520
rect 453946 488336 454002 488345
rect 453946 488271 454002 488280
rect 453960 487490 453988 488271
rect 453948 487484 454000 487490
rect 453948 487426 454000 487432
rect 453762 486976 453818 486985
rect 453762 486911 453818 486920
rect 453776 485858 453804 486911
rect 453764 485852 453816 485858
rect 453764 485794 453816 485800
rect 453946 485616 454002 485625
rect 453946 485551 454002 485560
rect 453960 484498 453988 485551
rect 453948 484492 454000 484498
rect 453948 484434 454000 484440
rect 453762 481536 453818 481545
rect 453762 481471 453818 481480
rect 453776 480282 453804 481471
rect 453764 480276 453816 480282
rect 453764 480218 453816 480224
rect 453762 478816 453818 478825
rect 453762 478751 453818 478760
rect 453776 477562 453804 478751
rect 453764 477556 453816 477562
rect 453764 477498 453816 477504
rect 453854 477456 453910 477465
rect 453854 477391 453910 477400
rect 453868 476134 453896 477391
rect 453856 476128 453908 476134
rect 453856 476070 453908 476076
rect 453946 476096 454002 476105
rect 453946 476031 454002 476040
rect 453960 474774 453988 476031
rect 453948 474768 454000 474774
rect 453948 474710 454000 474716
rect 453946 472696 454002 472705
rect 453946 472631 454002 472640
rect 453960 472394 453988 472631
rect 453948 472388 454000 472394
rect 453948 472330 454000 472336
rect 453762 471336 453818 471345
rect 453762 471271 453764 471280
rect 453816 471271 453818 471280
rect 453764 471242 453816 471248
rect 453946 469976 454002 469985
rect 453946 469911 454002 469920
rect 453960 469266 453988 469911
rect 453948 469260 454000 469266
rect 453948 469202 454000 469208
rect 453578 467256 453634 467265
rect 453578 467191 453634 467200
rect 453592 466682 453620 467191
rect 453580 466676 453632 466682
rect 453580 466618 453632 466624
rect 453946 463176 454002 463185
rect 453946 463111 454002 463120
rect 453960 462398 453988 463111
rect 453948 462392 454000 462398
rect 453948 462334 454000 462340
rect 453946 460456 454002 460465
rect 453946 460391 454002 460400
rect 453960 459610 453988 460391
rect 453948 459604 454000 459610
rect 453948 459546 454000 459552
rect 453670 456376 453726 456385
rect 453670 456311 453726 456320
rect 453684 455462 453712 456311
rect 453672 455456 453724 455462
rect 453672 455398 453724 455404
rect 453946 454336 454002 454345
rect 453946 454271 453948 454280
rect 454000 454271 454002 454280
rect 453948 454242 454000 454248
rect 453946 452976 454002 452985
rect 453946 452911 454002 452920
rect 453960 452674 453988 452911
rect 453948 452668 454000 452674
rect 453948 452610 454000 452616
rect 453578 450256 453634 450265
rect 453578 450191 453580 450200
rect 453632 450191 453634 450200
rect 453580 450162 453632 450168
rect 453946 444816 454002 444825
rect 453946 444751 453948 444760
rect 454000 444751 454002 444760
rect 453948 444722 454000 444728
rect 453946 440736 454002 440745
rect 453946 440671 454002 440680
rect 453960 440298 453988 440671
rect 453948 440292 454000 440298
rect 453948 440234 454000 440240
rect 453856 440224 453908 440230
rect 453856 440166 453908 440172
rect 453868 439385 453896 440166
rect 453854 439376 453910 439385
rect 453854 439311 453910 439320
rect 453946 438016 454002 438025
rect 453946 437951 454002 437960
rect 453960 437510 453988 437951
rect 453948 437504 454000 437510
rect 453948 437446 454000 437452
rect 453946 436656 454002 436665
rect 453946 436591 454002 436600
rect 453960 436150 453988 436591
rect 453948 436144 454000 436150
rect 453948 436086 454000 436092
rect 453670 435296 453726 435305
rect 453670 435231 453726 435240
rect 453684 435130 453712 435231
rect 453672 435124 453724 435130
rect 453672 435066 453724 435072
rect 453946 431896 454002 431905
rect 453946 431831 454002 431840
rect 453960 430642 453988 431831
rect 453948 430636 454000 430642
rect 453948 430578 454000 430584
rect 453946 429176 454002 429185
rect 453946 429111 454002 429120
rect 453960 427854 453988 429111
rect 453948 427848 454000 427854
rect 453948 427790 454000 427796
rect 453948 426488 454000 426494
rect 453946 426456 453948 426465
rect 454000 426456 454002 426465
rect 453946 426391 454002 426400
rect 453948 425128 454000 425134
rect 453946 425096 453948 425105
rect 454000 425096 454002 425105
rect 453946 425031 454002 425040
rect 453946 421016 454002 421025
rect 453946 420951 453948 420960
rect 454000 420951 454002 420960
rect 453948 420922 454000 420928
rect 453670 418296 453726 418305
rect 453670 418231 453672 418240
rect 453724 418231 453726 418240
rect 453672 418202 453724 418208
rect 453946 413536 454002 413545
rect 453946 413471 454002 413480
rect 453960 413234 453988 413471
rect 453948 413228 454000 413234
rect 453948 413170 454000 413176
rect 453762 408096 453818 408105
rect 453762 408031 453818 408040
rect 453776 407250 453804 408031
rect 453764 407244 453816 407250
rect 453764 407186 453816 407192
rect 453948 407108 454000 407114
rect 453948 407050 454000 407056
rect 453960 406745 453988 407050
rect 453946 406736 454002 406745
rect 453946 406671 454002 406680
rect 453762 405376 453818 405385
rect 453762 405311 453818 405320
rect 453776 404938 453804 405311
rect 453764 404932 453816 404938
rect 453764 404874 453816 404880
rect 453946 402656 454002 402665
rect 453946 402591 454002 402600
rect 453960 401674 453988 402591
rect 453948 401668 454000 401674
rect 453948 401610 454000 401616
rect 453762 399936 453818 399945
rect 453762 399871 453818 399880
rect 453776 398886 453804 399871
rect 453764 398880 453816 398886
rect 453764 398822 453816 398828
rect 453762 395856 453818 395865
rect 453762 395791 453818 395800
rect 453776 394738 453804 395791
rect 453764 394732 453816 394738
rect 453764 394674 453816 394680
rect 453762 394496 453818 394505
rect 453762 394431 453818 394440
rect 453776 393378 453804 394431
rect 453764 393372 453816 393378
rect 453764 393314 453816 393320
rect 453946 392456 454002 392465
rect 453946 392391 454002 392400
rect 453960 392018 453988 392391
rect 453948 392012 454000 392018
rect 453948 391954 454000 391960
rect 453946 389736 454002 389745
rect 453946 389671 454002 389680
rect 453960 389230 453988 389671
rect 453948 389224 454000 389230
rect 453948 389166 454000 389172
rect 453946 387016 454002 387025
rect 453946 386951 454002 386960
rect 453960 386714 453988 386951
rect 453948 386708 454000 386714
rect 453948 386650 454000 386656
rect 453948 385688 454000 385694
rect 453946 385656 453948 385665
rect 454000 385656 454002 385665
rect 453946 385591 454002 385600
rect 453946 384296 454002 384305
rect 453946 384231 454002 384240
rect 453960 383722 453988 384231
rect 453948 383716 454000 383722
rect 453948 383658 454000 383664
rect 453762 378856 453818 378865
rect 453762 378791 453764 378800
rect 453816 378791 453818 378800
rect 453764 378762 453816 378768
rect 453762 376136 453818 376145
rect 453762 376071 453818 376080
rect 453776 375970 453804 376071
rect 453764 375964 453816 375970
rect 453764 375906 453816 375912
rect 453946 372736 454002 372745
rect 453946 372671 453948 372680
rect 454000 372671 454002 372680
rect 453948 372642 454000 372648
rect 453762 371376 453818 371385
rect 453762 371311 453818 371320
rect 453776 371278 453804 371311
rect 453764 371272 453816 371278
rect 453764 371214 453816 371220
rect 453762 370016 453818 370025
rect 453762 369951 453818 369960
rect 453776 369918 453804 369951
rect 453764 369912 453816 369918
rect 453764 369854 453816 369860
rect 453762 368656 453818 368665
rect 453762 368591 453818 368600
rect 453776 368558 453804 368591
rect 453764 368552 453816 368558
rect 453764 368494 453816 368500
rect 453946 367296 454002 367305
rect 453946 367231 453948 367240
rect 454000 367231 454002 367240
rect 453948 367202 454000 367208
rect 453946 365936 454002 365945
rect 453946 365871 454002 365880
rect 453960 365770 453988 365871
rect 453948 365764 454000 365770
rect 453948 365706 454000 365712
rect 453762 364576 453818 364585
rect 453762 364511 453818 364520
rect 453776 364478 453804 364511
rect 453764 364472 453816 364478
rect 453764 364414 453816 364420
rect 453762 363216 453818 363225
rect 453762 363151 453818 363160
rect 453578 356416 453634 356425
rect 453578 356351 453634 356360
rect 453488 356040 453540 356046
rect 453488 355982 453540 355988
rect 453486 353696 453542 353705
rect 453486 353631 453542 353640
rect 453396 350396 453448 350402
rect 453396 350338 453448 350344
rect 453304 347744 453356 347750
rect 453304 347686 453356 347692
rect 453210 346216 453266 346225
rect 453210 346151 453266 346160
rect 453224 319462 453252 346151
rect 453500 334626 453528 353631
rect 453592 338337 453620 356351
rect 453670 350296 453726 350305
rect 453670 350231 453726 350240
rect 453578 338328 453634 338337
rect 453578 338263 453634 338272
rect 453488 334620 453540 334626
rect 453488 334562 453540 334568
rect 453212 319456 453264 319462
rect 453212 319398 453264 319404
rect 453120 308440 453172 308446
rect 453120 308382 453172 308388
rect 452844 180124 452896 180130
rect 452844 180066 452896 180072
rect 452752 87644 452804 87650
rect 452752 87586 452804 87592
rect 453684 35222 453712 350231
rect 453776 326466 453804 363151
rect 453946 361856 454002 361865
rect 453946 361791 454002 361800
rect 453960 361622 453988 361791
rect 453948 361616 454000 361622
rect 453948 361558 454000 361564
rect 453946 359136 454002 359145
rect 453946 359071 454002 359080
rect 453960 358834 453988 359071
rect 453948 358828 454000 358834
rect 453948 358770 454000 358776
rect 453946 357776 454002 357785
rect 453946 357711 454002 357720
rect 453960 357542 453988 357711
rect 453948 357536 454000 357542
rect 453948 357478 454000 357484
rect 453946 348936 454002 348945
rect 453946 348871 454002 348880
rect 453960 347818 453988 348871
rect 454052 348838 454080 554746
rect 455696 549500 455748 549506
rect 455696 549442 455748 549448
rect 455604 544060 455656 544066
rect 455604 544002 455656 544008
rect 454130 526416 454186 526425
rect 454130 526351 454186 526360
rect 454040 348832 454092 348838
rect 454040 348774 454092 348780
rect 453948 347812 454000 347818
rect 453948 347754 454000 347760
rect 454040 347744 454092 347750
rect 454040 347686 454092 347692
rect 453948 347608 454000 347614
rect 453946 347576 453948 347585
rect 454000 347576 454002 347585
rect 453946 347511 454002 347520
rect 453946 343496 454002 343505
rect 453946 343431 454002 343440
rect 453960 342310 453988 343431
rect 453948 342304 454000 342310
rect 453948 342246 454000 342252
rect 453946 342136 454002 342145
rect 453946 342071 453948 342080
rect 454000 342071 454002 342080
rect 453948 342042 454000 342048
rect 454052 341465 454080 347686
rect 454038 341456 454094 341465
rect 454038 341391 454094 341400
rect 454144 337618 454172 526351
rect 454408 468580 454460 468586
rect 454408 468522 454460 468528
rect 454222 465896 454278 465905
rect 454222 465831 454278 465840
rect 454132 337612 454184 337618
rect 454132 337554 454184 337560
rect 453764 326460 453816 326466
rect 453764 326402 453816 326408
rect 454236 323610 454264 465831
rect 454316 458448 454368 458454
rect 454316 458390 454368 458396
rect 454224 323604 454276 323610
rect 454224 323546 454276 323552
rect 454328 318102 454356 458390
rect 454420 327758 454448 468522
rect 455420 464228 455472 464234
rect 455420 464170 455472 464176
rect 454500 447500 454552 447506
rect 454500 447442 454552 447448
rect 454512 330682 454540 447442
rect 454592 408876 454644 408882
rect 454592 408818 454644 408824
rect 454604 336326 454632 408818
rect 454684 400240 454736 400246
rect 454684 400182 454736 400188
rect 454696 337414 454724 400182
rect 454960 350396 455012 350402
rect 454960 350338 455012 350344
rect 454868 343936 454920 343942
rect 454868 343878 454920 343884
rect 454684 337408 454736 337414
rect 454684 337350 454736 337356
rect 454592 336320 454644 336326
rect 454592 336262 454644 336268
rect 454500 330676 454552 330682
rect 454500 330618 454552 330624
rect 454408 327752 454460 327758
rect 454408 327694 454460 327700
rect 454316 318096 454368 318102
rect 454316 318038 454368 318044
rect 453672 35216 453724 35222
rect 453672 35158 453724 35164
rect 454880 6914 454908 343878
rect 454972 342378 455000 350338
rect 454960 342372 455012 342378
rect 454960 342314 455012 342320
rect 455432 47598 455460 464170
rect 455512 416900 455564 416906
rect 455512 416842 455564 416848
rect 455524 174554 455552 416842
rect 455616 327826 455644 544002
rect 455708 337210 455736 549442
rect 455788 524748 455840 524754
rect 455788 524690 455840 524696
rect 455696 337204 455748 337210
rect 455696 337146 455748 337152
rect 455800 330614 455828 524690
rect 455972 466676 456024 466682
rect 455972 466618 456024 466624
rect 455880 450220 455932 450226
rect 455880 450162 455932 450168
rect 455788 330608 455840 330614
rect 455788 330550 455840 330556
rect 455604 327820 455656 327826
rect 455604 327762 455656 327768
rect 455892 297430 455920 450162
rect 455984 334966 456012 466618
rect 456064 435124 456116 435130
rect 456064 435066 456116 435072
rect 455972 334960 456024 334966
rect 455972 334902 456024 334908
rect 456076 307086 456104 435066
rect 456156 418260 456208 418266
rect 456156 418202 456208 418208
rect 456168 326398 456196 418202
rect 456248 407244 456300 407250
rect 456248 407186 456300 407192
rect 456260 331974 456288 407186
rect 456800 357536 456852 357542
rect 456800 357478 456852 357484
rect 456812 337754 456840 357478
rect 456800 337748 456852 337754
rect 456800 337690 456852 337696
rect 456904 335646 456932 559302
rect 456996 385694 457024 562294
rect 459008 559496 459060 559502
rect 459008 559438 459060 559444
rect 457076 559428 457128 559434
rect 457076 559370 457128 559376
rect 456984 385688 457036 385694
rect 456984 385630 457036 385636
rect 456984 372700 457036 372706
rect 456984 372642 457036 372648
rect 456892 335640 456944 335646
rect 456892 335582 456944 335588
rect 456248 331968 456300 331974
rect 456248 331910 456300 331916
rect 456156 326392 456208 326398
rect 456156 326334 456208 326340
rect 456064 307080 456116 307086
rect 456064 307022 456116 307028
rect 456798 300112 456854 300121
rect 456798 300047 456854 300056
rect 455880 297424 455932 297430
rect 455880 297366 455932 297372
rect 455512 174548 455564 174554
rect 455512 174490 455564 174496
rect 455420 47592 455472 47598
rect 455420 47534 455472 47540
rect 454512 6886 454908 6914
rect 453304 3596 453356 3602
rect 453304 3538 453356 3544
rect 452384 3324 452436 3330
rect 452384 3266 452436 3272
rect 451924 3120 451976 3126
rect 451924 3062 451976 3068
rect 453316 480 453344 3538
rect 453580 3528 453632 3534
rect 453580 3470 453632 3476
rect 453592 3330 453620 3470
rect 453580 3324 453632 3330
rect 453580 3266 453632 3272
rect 454512 480 454540 6886
rect 455696 3732 455748 3738
rect 455696 3674 455748 3680
rect 455708 480 455736 3674
rect 456812 3346 456840 300047
rect 456890 261488 456946 261497
rect 456890 261423 456946 261432
rect 456904 3534 456932 261423
rect 456996 33114 457024 372642
rect 457088 338881 457116 559370
rect 458364 559224 458416 559230
rect 458364 559166 458416 559172
rect 457628 546576 457680 546582
rect 457628 546518 457680 546524
rect 457168 520940 457220 520946
rect 457168 520882 457220 520888
rect 457074 338872 457130 338881
rect 457074 338807 457130 338816
rect 457180 322318 457208 520882
rect 457260 498500 457312 498506
rect 457260 498442 457312 498448
rect 457272 336054 457300 498442
rect 457352 454300 457404 454306
rect 457352 454242 457404 454248
rect 457260 336048 457312 336054
rect 457260 335990 457312 335996
rect 457364 324970 457392 454242
rect 457444 386708 457496 386714
rect 457444 386650 457496 386656
rect 457456 333402 457484 386650
rect 457536 378820 457588 378826
rect 457536 378762 457588 378768
rect 457548 339289 457576 378762
rect 457534 339280 457590 339289
rect 457534 339215 457590 339224
rect 457444 333396 457496 333402
rect 457444 333338 457496 333344
rect 457352 324964 457404 324970
rect 457352 324906 457404 324912
rect 457168 322312 457220 322318
rect 457168 322254 457220 322260
rect 457640 309806 457668 546518
rect 458272 471300 458324 471306
rect 458272 471242 458324 471248
rect 458180 342100 458232 342106
rect 458180 342042 458232 342048
rect 458192 333266 458220 342042
rect 458180 333260 458232 333266
rect 458180 333202 458232 333208
rect 457628 309800 457680 309806
rect 457628 309742 457680 309748
rect 458284 239426 458312 471242
rect 458376 339697 458404 559166
rect 458456 487484 458508 487490
rect 458456 487426 458508 487432
rect 458362 339688 458418 339697
rect 458362 339623 458418 339632
rect 458468 294642 458496 487426
rect 458548 484492 458600 484498
rect 458548 484434 458600 484440
rect 458560 302938 458588 484434
rect 458640 472388 458692 472394
rect 458640 472330 458692 472336
rect 458652 312594 458680 472330
rect 458732 413228 458784 413234
rect 458732 413170 458784 413176
rect 458744 337686 458772 413170
rect 458824 375964 458876 375970
rect 458824 375906 458876 375912
rect 458836 338609 458864 375906
rect 458916 367260 458968 367266
rect 458916 367202 458968 367208
rect 458822 338600 458878 338609
rect 458822 338535 458878 338544
rect 458732 337680 458784 337686
rect 458732 337622 458784 337628
rect 458928 333441 458956 367202
rect 458914 333432 458970 333441
rect 458914 333367 458970 333376
rect 458640 312588 458692 312594
rect 458640 312530 458692 312536
rect 458548 302932 458600 302938
rect 458548 302874 458600 302880
rect 458456 294636 458508 294642
rect 458456 294578 458508 294584
rect 458272 239420 458324 239426
rect 458272 239362 458324 239368
rect 456984 33108 457036 33114
rect 456984 33050 457036 33056
rect 456892 3528 456944 3534
rect 456892 3470 456944 3476
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 456812 3318 456932 3346
rect 456904 480 456932 3318
rect 458100 480 458128 3470
rect 459020 3330 459048 559438
rect 459560 556640 459612 556646
rect 459560 556582 459612 556588
rect 459572 4078 459600 556582
rect 459664 347614 459692 700470
rect 462332 699718 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 461676 699712 461728 699718
rect 461676 699654 461728 699660
rect 462320 699712 462372 699718
rect 462320 699654 462372 699660
rect 459928 559700 459980 559706
rect 459928 559642 459980 559648
rect 459836 482792 459888 482798
rect 459836 482734 459888 482740
rect 459744 356040 459796 356046
rect 459744 355982 459796 355988
rect 459652 347608 459704 347614
rect 459652 347550 459704 347556
rect 459652 39364 459704 39370
rect 459652 39306 459704 39312
rect 459560 4072 459612 4078
rect 459560 4014 459612 4020
rect 459192 3868 459244 3874
rect 459192 3810 459244 3816
rect 459008 3324 459060 3330
rect 459008 3266 459060 3272
rect 459204 480 459232 3810
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459664 354 459692 39306
rect 459756 3806 459784 355982
rect 459848 255270 459876 482734
rect 459940 336190 459968 559642
rect 461400 559632 461452 559638
rect 461400 559574 461452 559580
rect 460940 559564 460992 559570
rect 460940 559506 460992 559512
rect 460204 558136 460256 558142
rect 460204 558078 460256 558084
rect 460020 444780 460072 444786
rect 460020 444722 460072 444728
rect 460032 336394 460060 444722
rect 460112 404932 460164 404938
rect 460112 404874 460164 404880
rect 460020 336388 460072 336394
rect 460020 336330 460072 336336
rect 459928 336184 459980 336190
rect 459928 336126 459980 336132
rect 460124 336025 460152 404874
rect 460110 336016 460166 336025
rect 460110 335951 460166 335960
rect 459836 255264 459888 255270
rect 459836 255206 459888 255212
rect 459744 3800 459796 3806
rect 459744 3742 459796 3748
rect 460216 3534 460244 558078
rect 460388 382900 460440 382906
rect 460388 382842 460440 382848
rect 460296 378208 460348 378214
rect 460296 378150 460348 378156
rect 460308 333674 460336 378150
rect 460400 338745 460428 382842
rect 460386 338736 460442 338745
rect 460386 338671 460442 338680
rect 460296 333668 460348 333674
rect 460296 333610 460348 333616
rect 460952 3670 460980 559506
rect 461124 556776 461176 556782
rect 461124 556718 461176 556724
rect 461032 556436 461084 556442
rect 461032 556378 461084 556384
rect 461044 4010 461072 556378
rect 461032 4004 461084 4010
rect 461032 3946 461084 3952
rect 460940 3664 460992 3670
rect 460940 3606 460992 3612
rect 461136 3602 461164 556718
rect 461216 532772 461268 532778
rect 461216 532714 461268 532720
rect 461228 293962 461256 532714
rect 461308 436144 461360 436150
rect 461308 436086 461360 436092
rect 461216 293956 461268 293962
rect 461216 293898 461268 293904
rect 461320 202842 461348 436086
rect 461412 336530 461440 559574
rect 461584 521688 461636 521694
rect 461584 521630 461636 521636
rect 461492 394732 461544 394738
rect 461492 394674 461544 394680
rect 461400 336524 461452 336530
rect 461400 336466 461452 336472
rect 461504 267714 461532 394674
rect 461492 267708 461544 267714
rect 461492 267650 461544 267656
rect 461308 202836 461360 202842
rect 461308 202778 461360 202784
rect 461596 6866 461624 521630
rect 461688 339017 461716 699654
rect 465724 696992 465776 696998
rect 465724 696934 465776 696940
rect 464528 560788 464580 560794
rect 464528 560730 464580 560736
rect 463790 559328 463846 559337
rect 463790 559263 463846 559272
rect 462412 559020 462464 559026
rect 462412 558962 462464 558968
rect 461768 364404 461820 364410
rect 461768 364346 461820 364352
rect 461674 339008 461730 339017
rect 461674 338943 461730 338952
rect 461780 336666 461808 364346
rect 462320 361616 462372 361622
rect 462320 361558 462372 361564
rect 461768 336660 461820 336666
rect 461768 336602 461820 336608
rect 462332 333334 462360 361558
rect 462320 333328 462372 333334
rect 462320 333270 462372 333276
rect 461676 9036 461728 9042
rect 461676 8978 461728 8984
rect 461584 6860 461636 6866
rect 461584 6802 461636 6808
rect 461124 3596 461176 3602
rect 461124 3538 461176 3544
rect 460204 3528 460256 3534
rect 461688 3482 461716 8978
rect 462424 4146 462452 558962
rect 462504 556844 462556 556850
rect 462504 556786 462556 556792
rect 462412 4140 462464 4146
rect 462412 4082 462464 4088
rect 460204 3470 460256 3476
rect 461596 3454 461716 3482
rect 461596 480 461624 3454
rect 462516 3398 462544 556786
rect 462596 556708 462648 556714
rect 462596 556650 462648 556656
rect 462608 3738 462636 556650
rect 462688 541000 462740 541006
rect 462688 540942 462740 540948
rect 462700 333810 462728 540942
rect 463148 536852 463200 536858
rect 463148 536794 463200 536800
rect 462780 509312 462832 509318
rect 462780 509254 462832 509260
rect 462792 337822 462820 509254
rect 462872 455456 462924 455462
rect 462872 455398 462924 455404
rect 462780 337816 462832 337822
rect 462780 337758 462832 337764
rect 462884 337278 462912 455398
rect 462964 429888 463016 429894
rect 462964 429830 463016 429836
rect 462872 337272 462924 337278
rect 462872 337214 462924 337220
rect 462976 336462 463004 429830
rect 463056 401668 463108 401674
rect 463056 401610 463108 401616
rect 462964 336456 463016 336462
rect 462964 336398 463016 336404
rect 463068 336258 463096 401610
rect 463056 336252 463108 336258
rect 463056 336194 463108 336200
rect 462688 333804 462740 333810
rect 462688 333746 462740 333752
rect 463160 6914 463188 536794
rect 463700 364472 463752 364478
rect 463700 364414 463752 364420
rect 463712 333198 463740 364414
rect 463700 333192 463752 333198
rect 463700 333134 463752 333140
rect 462792 6886 463188 6914
rect 462596 3732 462648 3738
rect 462596 3674 462648 3680
rect 462504 3392 462556 3398
rect 462504 3334 462556 3340
rect 462792 480 462820 6886
rect 463804 3233 463832 559263
rect 463974 559192 464030 559201
rect 463974 559127 464030 559136
rect 463884 420980 463936 420986
rect 463884 420922 463936 420928
rect 463896 3942 463924 420922
rect 463988 337521 464016 559127
rect 464068 559088 464120 559094
rect 464068 559030 464120 559036
rect 464080 337890 464108 559030
rect 464252 503736 464304 503742
rect 464252 503678 464304 503684
rect 464160 365764 464212 365770
rect 464160 365706 464212 365712
rect 464068 337884 464120 337890
rect 464068 337826 464120 337832
rect 463974 337512 464030 337521
rect 463974 337447 464030 337456
rect 464172 189038 464200 365706
rect 464264 337142 464292 503678
rect 464344 488572 464396 488578
rect 464344 488514 464396 488520
rect 464252 337136 464304 337142
rect 464252 337078 464304 337084
rect 464160 189032 464212 189038
rect 464160 188974 464212 188980
rect 463976 18624 464028 18630
rect 463976 18566 464028 18572
rect 463884 3936 463936 3942
rect 463884 3878 463936 3884
rect 463790 3224 463846 3233
rect 463790 3159 463846 3168
rect 463988 480 464016 18566
rect 464356 9654 464384 488514
rect 464436 393372 464488 393378
rect 464436 393314 464488 393320
rect 464448 336598 464476 393314
rect 464436 336592 464488 336598
rect 464436 336534 464488 336540
rect 464344 9648 464396 9654
rect 464344 9590 464396 9596
rect 464540 3194 464568 560730
rect 465262 559464 465318 559473
rect 465262 559399 465318 559408
rect 465172 557796 465224 557802
rect 465172 557738 465224 557744
rect 465184 16574 465212 557738
rect 465276 333470 465304 559399
rect 465356 559292 465408 559298
rect 465356 559234 465408 559240
rect 465368 337346 465396 559234
rect 465736 513330 465764 696934
rect 465816 560856 465868 560862
rect 465816 560798 465868 560804
rect 465724 513324 465776 513330
rect 465724 513266 465776 513272
rect 465724 477556 465776 477562
rect 465724 477498 465776 477504
rect 465448 452668 465500 452674
rect 465448 452610 465500 452616
rect 465356 337340 465408 337346
rect 465356 337282 465408 337288
rect 465460 336433 465488 452610
rect 465540 398880 465592 398886
rect 465540 398822 465592 398828
rect 465446 336424 465502 336433
rect 465446 336359 465502 336368
rect 465264 333464 465316 333470
rect 465264 333406 465316 333412
rect 465552 333305 465580 398822
rect 465632 389224 465684 389230
rect 465632 389166 465684 389172
rect 465644 338230 465672 389166
rect 465632 338224 465684 338230
rect 465632 338166 465684 338172
rect 465538 333296 465594 333305
rect 465538 333231 465594 333240
rect 465262 36544 465318 36553
rect 465262 36479 465318 36488
rect 465092 16546 465212 16574
rect 465092 3262 465120 16546
rect 465172 9648 465224 9654
rect 465172 9590 465224 9596
rect 465080 3256 465132 3262
rect 465080 3198 465132 3204
rect 464528 3188 464580 3194
rect 464528 3130 464580 3136
rect 465184 480 465212 9590
rect 465276 6914 465304 36479
rect 465736 14482 465764 477498
rect 465828 16574 465856 560798
rect 474002 559600 474058 559609
rect 474002 559535 474058 559544
rect 469864 558952 469916 558958
rect 469864 558894 469916 558900
rect 466460 557932 466512 557938
rect 466460 557874 466512 557880
rect 466472 16574 466500 557874
rect 469220 556980 469272 556986
rect 469220 556922 469272 556928
rect 468576 553444 468628 553450
rect 468576 553386 468628 553392
rect 468484 542428 468536 542434
rect 468484 542370 468536 542376
rect 467840 268456 467892 268462
rect 467840 268398 467892 268404
rect 467852 16574 467880 268398
rect 465828 16546 465948 16574
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 465724 14476 465776 14482
rect 465724 14418 465776 14424
rect 465276 6886 465856 6914
rect 460358 354 460470 480
rect 459664 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 6886
rect 465920 3641 465948 16546
rect 465906 3632 465962 3641
rect 465906 3567 465962 3576
rect 467484 480 467512 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 468496 8974 468524 542370
rect 468588 299470 468616 553386
rect 468576 299464 468628 299470
rect 468576 299406 468628 299412
rect 469232 16574 469260 556922
rect 469876 138718 469904 558894
rect 472624 558068 472676 558074
rect 472624 558010 472676 558016
rect 471980 527196 472032 527202
rect 471980 527138 472032 527144
rect 471336 484424 471388 484430
rect 471336 484366 471388 484372
rect 471244 342304 471296 342310
rect 471244 342246 471296 342252
rect 469864 138712 469916 138718
rect 469864 138654 469916 138660
rect 470600 43444 470652 43450
rect 470600 43386 470652 43392
rect 469232 16546 469904 16574
rect 468484 8968 468536 8974
rect 468484 8910 468536 8916
rect 469876 480 469904 16546
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 43386
rect 471256 3602 471284 342246
rect 471348 333878 471376 484366
rect 471336 333872 471388 333878
rect 471336 333814 471388 333820
rect 471992 16574 472020 527138
rect 471992 16546 472296 16574
rect 471244 3596 471296 3602
rect 471244 3538 471296 3544
rect 472268 480 472296 16546
rect 472636 3058 472664 558010
rect 474016 33114 474044 559535
rect 475476 518968 475528 518974
rect 475476 518910 475528 518916
rect 475384 462392 475436 462398
rect 475384 462334 475436 462340
rect 474740 91792 474792 91798
rect 474740 91734 474792 91740
rect 474004 33108 474056 33114
rect 474004 33050 474056 33056
rect 473452 22772 473504 22778
rect 473452 22714 473504 22720
rect 472624 3052 472676 3058
rect 472624 2994 472676 3000
rect 473464 480 473492 22714
rect 474752 16574 474780 91734
rect 474752 16546 475332 16574
rect 475304 3482 475332 16546
rect 475396 4146 475424 462334
rect 475488 193186 475516 518910
rect 476764 371272 476816 371278
rect 476764 371214 476816 371220
rect 475476 193180 475528 193186
rect 475476 193122 475528 193128
rect 476118 37904 476174 37913
rect 476118 37839 476174 37848
rect 476132 16574 476160 37839
rect 476132 16546 476528 16574
rect 475384 4140 475436 4146
rect 475384 4082 475436 4088
rect 475936 4140 475988 4146
rect 475936 4082 475988 4088
rect 475304 3454 475792 3482
rect 474556 3052 474608 3058
rect 474556 2994 474608 3000
rect 474568 480 474596 2994
rect 475764 480 475792 3454
rect 475948 3330 475976 4082
rect 475936 3324 475988 3330
rect 475936 3266 475988 3272
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 476776 4826 476804 371214
rect 477512 333742 477540 702406
rect 485044 590708 485096 590714
rect 485044 590650 485096 590656
rect 483020 560924 483072 560930
rect 483020 560866 483072 560872
rect 480260 560652 480312 560658
rect 480260 560594 480312 560600
rect 479524 536852 479576 536858
rect 479524 536794 479576 536800
rect 478880 347812 478932 347818
rect 478880 347754 478932 347760
rect 477500 333736 477552 333742
rect 477500 333678 477552 333684
rect 477500 325100 477552 325106
rect 477500 325042 477552 325048
rect 477512 16574 477540 325042
rect 477512 16546 478184 16574
rect 476764 4820 476816 4826
rect 476764 4762 476816 4768
rect 478156 480 478184 16546
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 347754
rect 479536 333606 479564 536794
rect 479524 333600 479576 333606
rect 479524 333542 479576 333548
rect 480272 16574 480300 560594
rect 481732 558204 481784 558210
rect 481732 558146 481784 558152
rect 480904 485852 480956 485858
rect 480904 485794 480956 485800
rect 480916 100706 480944 485794
rect 480904 100700 480956 100706
rect 480904 100642 480956 100648
rect 481744 16574 481772 558146
rect 483032 16574 483060 560866
rect 485056 336734 485084 590650
rect 494072 562426 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700330 527220 703520
rect 543476 700466 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 498844 683188 498896 683194
rect 498844 683130 498896 683136
rect 494060 562420 494112 562426
rect 494060 562362 494112 562368
rect 487160 560584 487212 560590
rect 487160 560526 487212 560532
rect 486516 470620 486568 470626
rect 486516 470562 486568 470568
rect 486424 368552 486476 368558
rect 486424 368494 486476 368500
rect 485044 336728 485096 336734
rect 485044 336670 485096 336676
rect 484400 295996 484452 296002
rect 484400 295938 484452 295944
rect 484412 16574 484440 295938
rect 486436 16574 486464 368494
rect 486528 336122 486556 470562
rect 486516 336116 486568 336122
rect 486516 336058 486568 336064
rect 480272 16546 480576 16574
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 486436 16546 486556 16574
rect 480548 480 480576 16546
rect 481732 3324 481784 3330
rect 481732 3266 481784 3272
rect 481744 480 481772 3266
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486528 3602 486556 16546
rect 486424 3596 486476 3602
rect 486424 3538 486476 3544
rect 486516 3596 486568 3602
rect 486516 3538 486568 3544
rect 486436 480 486464 3538
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 560526
rect 492680 557728 492732 557734
rect 492680 557670 492732 557676
rect 489184 437504 489236 437510
rect 489184 437446 489236 437452
rect 489196 31074 489224 437446
rect 491944 418192 491996 418198
rect 491944 418134 491996 418140
rect 491956 407114 491984 418134
rect 491944 407108 491996 407114
rect 491944 407050 491996 407056
rect 491300 392012 491352 392018
rect 491300 391954 491352 391960
rect 489920 46232 489972 46238
rect 489920 46174 489972 46180
rect 489184 31068 489236 31074
rect 489184 31010 489236 31016
rect 488540 29640 488592 29646
rect 488540 29582 488592 29588
rect 488552 16574 488580 29582
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 480 489960 46174
rect 491312 16574 491340 391954
rect 492692 16574 492720 557670
rect 496820 557660 496872 557666
rect 496820 557602 496872 557608
rect 495440 556912 495492 556918
rect 495440 556854 495492 556860
rect 494060 426488 494112 426494
rect 494060 426430 494112 426436
rect 494072 16574 494100 426430
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 491116 8968 491168 8974
rect 491116 8910 491168 8916
rect 491128 480 491156 8910
rect 492324 480 492352 16546
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 556854
rect 496832 16574 496860 557602
rect 498856 492658 498884 683130
rect 502984 643136 503036 643142
rect 502984 643078 503036 643084
rect 500960 562148 501012 562154
rect 500960 562090 501012 562096
rect 500224 514820 500276 514826
rect 500224 514762 500276 514768
rect 498844 492652 498896 492658
rect 498844 492594 498896 492600
rect 498200 305652 498252 305658
rect 498200 305594 498252 305600
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 305594
rect 499396 4820 499448 4826
rect 499396 4762 499448 4768
rect 499408 480 499436 4762
rect 500236 3738 500264 514762
rect 500972 16574 501000 562090
rect 502996 440230 503024 643078
rect 531412 562080 531464 562086
rect 531412 562022 531464 562028
rect 507124 560448 507176 560454
rect 507124 560390 507176 560396
rect 503720 558000 503772 558006
rect 503720 557942 503772 557948
rect 502984 440224 503036 440230
rect 502984 440166 503036 440172
rect 502984 383716 503036 383722
rect 502984 383658 503036 383664
rect 502340 294704 502392 294710
rect 502340 294646 502392 294652
rect 500972 16546 501368 16574
rect 500224 3732 500276 3738
rect 500224 3674 500276 3680
rect 500592 3596 500644 3602
rect 500592 3538 500644 3544
rect 500604 480 500632 3538
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502352 6914 502380 294646
rect 502996 8974 503024 383658
rect 502984 8968 503036 8974
rect 502984 8910 503036 8916
rect 502352 6886 503024 6914
rect 502996 480 503024 6886
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 557942
rect 504364 459604 504416 459610
rect 504364 459546 504416 459552
rect 504376 3670 504404 459546
rect 505098 331800 505154 331809
rect 505098 331735 505154 331744
rect 505112 16574 505140 331735
rect 507136 46918 507164 560390
rect 527824 560380 527876 560386
rect 527824 560322 527876 560328
rect 524420 557864 524472 557870
rect 524420 557806 524472 557812
rect 518900 556504 518952 556510
rect 518900 556446 518952 556452
rect 512000 556368 512052 556374
rect 512000 556310 512052 556316
rect 507858 329216 507914 329225
rect 507858 329151 507914 329160
rect 507124 46912 507176 46918
rect 507124 46854 507176 46860
rect 506480 31068 506532 31074
rect 506480 31010 506532 31016
rect 505112 16546 505416 16574
rect 504364 3664 504416 3670
rect 504364 3606 504416 3612
rect 505388 480 505416 16546
rect 506492 480 506520 31010
rect 507872 16574 507900 329151
rect 510620 320884 510672 320890
rect 510620 320826 510672 320832
rect 510632 16574 510660 320826
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 507676 7812 507728 7818
rect 507676 7754 507728 7760
rect 507688 480 507716 7754
rect 508884 480 508912 16546
rect 509608 14476 509660 14482
rect 509608 14418 509660 14424
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509620 354 509648 14418
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 556310
rect 513380 556300 513432 556306
rect 513380 556242 513432 556248
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 556242
rect 517518 329080 517574 329089
rect 517518 329015 517574 329024
rect 516140 290488 516192 290494
rect 516140 290430 516192 290436
rect 514760 24132 514812 24138
rect 514760 24074 514812 24080
rect 514772 480 514800 24074
rect 516152 16574 516180 290430
rect 517532 16574 517560 329015
rect 518912 16574 518940 556446
rect 520924 535492 520976 535498
rect 520924 535434 520976 535440
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 515496 10328 515548 10334
rect 515496 10270 515548 10276
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 354 515536 10270
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 520740 8968 520792 8974
rect 520740 8910 520792 8916
rect 520752 480 520780 8910
rect 520936 3602 520964 535434
rect 523130 316840 523186 316849
rect 523130 316775 523186 316784
rect 521658 170368 521714 170377
rect 521658 170303 521714 170312
rect 520924 3596 520976 3602
rect 520924 3538 520976 3544
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521672 354 521700 170303
rect 523144 16574 523172 316775
rect 524432 16574 524460 557806
rect 526444 430636 526496 430642
rect 526444 430578 526496 430584
rect 525064 427848 525116 427854
rect 525064 427790 525116 427796
rect 523144 16546 523816 16574
rect 524432 16546 525012 16574
rect 523040 3460 523092 3466
rect 523040 3402 523092 3408
rect 523052 480 523080 3402
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 524984 3482 525012 16546
rect 525076 3806 525104 427790
rect 526168 11756 526220 11762
rect 526168 11698 526220 11704
rect 525064 3800 525116 3806
rect 525064 3742 525116 3748
rect 524984 3454 525472 3482
rect 525444 480 525472 3454
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 11698
rect 526456 8974 526484 430578
rect 527836 153202 527864 560322
rect 529204 469260 529256 469266
rect 529204 469202 529256 469208
rect 527824 153196 527876 153202
rect 527824 153138 527876 153144
rect 527180 152516 527232 152522
rect 527180 152458 527232 152464
rect 527192 16574 527220 152458
rect 528560 47660 528612 47666
rect 528560 47602 528612 47608
rect 527192 16546 527864 16574
rect 526444 8968 526496 8974
rect 526444 8910 526496 8916
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 47602
rect 529216 3466 529244 469202
rect 531424 6914 531452 562022
rect 540980 562012 541032 562018
rect 540980 561954 541032 561960
rect 538864 560516 538916 560522
rect 538864 560458 538916 560464
rect 536840 545148 536892 545154
rect 536840 545090 536892 545096
rect 534080 369912 534132 369918
rect 534080 369854 534132 369860
rect 533344 303000 533396 303006
rect 533344 302942 533396 302948
rect 533252 15904 533304 15910
rect 533252 15846 533304 15852
rect 531332 6886 531452 6914
rect 530122 3768 530178 3777
rect 530122 3703 530178 3712
rect 529204 3460 529256 3466
rect 529204 3402 529256 3408
rect 530136 480 530164 3703
rect 531332 480 531360 6886
rect 532516 3732 532568 3738
rect 532516 3674 532568 3680
rect 532528 480 532556 3674
rect 533264 3482 533292 15846
rect 533356 3738 533384 302942
rect 534092 16574 534120 369854
rect 536852 16574 536880 545090
rect 538220 25560 538272 25566
rect 538220 25502 538272 25508
rect 534092 16546 534488 16574
rect 536852 16546 537248 16574
rect 533344 3732 533396 3738
rect 533344 3674 533396 3680
rect 533264 3454 533752 3482
rect 533724 480 533752 3454
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536104 3732 536156 3738
rect 536104 3674 536156 3680
rect 536116 480 536144 3674
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 25502
rect 538876 20670 538904 560458
rect 538864 20664 538916 20670
rect 538864 20606 538916 20612
rect 540992 16574 541020 561954
rect 558932 560998 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580354 577688 580410 577697
rect 580354 577623 580410 577632
rect 580368 570654 580396 577623
rect 580356 570648 580408 570654
rect 580356 570590 580408 570596
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 572812 561944 572864 561950
rect 572812 561886 572864 561892
rect 569960 561740 570012 561746
rect 569960 561682 570012 561688
rect 558920 560992 558972 560998
rect 558920 560934 558972 560940
rect 565820 557592 565872 557598
rect 560298 557560 560354 557569
rect 565820 557534 565872 557540
rect 560298 557495 560354 557504
rect 557538 556472 557594 556481
rect 557538 556407 557594 556416
rect 550638 556336 550694 556345
rect 550638 556271 550694 556280
rect 541624 510672 541676 510678
rect 541624 510614 541676 510620
rect 541636 425066 541664 510614
rect 548524 499588 548576 499594
rect 548524 499530 548576 499536
rect 543004 480276 543056 480282
rect 543004 480218 543056 480224
rect 541624 425060 541676 425066
rect 541624 425002 541676 425008
rect 540992 16546 542032 16574
rect 540796 8968 540848 8974
rect 540796 8910 540848 8916
rect 539600 3664 539652 3670
rect 539600 3606 539652 3612
rect 539612 480 539640 3606
rect 540808 480 540836 8910
rect 542004 480 542032 16546
rect 543016 6934 543044 480218
rect 544384 440292 544436 440298
rect 544384 440234 544436 440240
rect 544396 16574 544424 440234
rect 547880 305720 547932 305726
rect 547880 305662 547932 305668
rect 547892 16574 547920 305662
rect 544396 16546 544516 16574
rect 547892 16546 548472 16574
rect 544384 13116 544436 13122
rect 544384 13058 544436 13064
rect 543188 7676 543240 7682
rect 543188 7618 543240 7624
rect 543004 6928 543056 6934
rect 543004 6870 543056 6876
rect 543200 480 543228 7618
rect 544396 480 544424 13058
rect 544488 4214 544516 16546
rect 547880 6928 547932 6934
rect 547880 6870 547932 6876
rect 544476 4208 544528 4214
rect 544476 4150 544528 4156
rect 545488 4208 545540 4214
rect 545488 4150 545540 4156
rect 545500 480 545528 4150
rect 546684 3528 546736 3534
rect 546684 3470 546736 3476
rect 546696 480 546724 3470
rect 547892 480 547920 6870
rect 548444 490 548472 16546
rect 548536 3058 548564 499530
rect 549904 476128 549956 476134
rect 549904 476070 549956 476076
rect 549260 284980 549312 284986
rect 549260 284922 549312 284928
rect 549272 6914 549300 284922
rect 549916 7614 549944 476070
rect 550652 16574 550680 556271
rect 556804 474768 556856 474774
rect 556804 474710 556856 474716
rect 555424 425128 555476 425134
rect 555424 425070 555476 425076
rect 552018 318200 552074 318209
rect 552018 318135 552074 318144
rect 552032 16574 552060 318135
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 549904 7608 549956 7614
rect 549904 7550 549956 7556
rect 549272 6886 550312 6914
rect 548524 3052 548576 3058
rect 548524 2994 548576 3000
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548444 462 548656 490
rect 550284 480 550312 6886
rect 548628 354 548656 462
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553766 6216 553822 6225
rect 553766 6151 553822 6160
rect 553780 480 553808 6151
rect 555436 3670 555464 425070
rect 556816 313274 556844 474710
rect 556804 313268 556856 313274
rect 556804 313210 556856 313216
rect 556252 291848 556304 291854
rect 556252 291790 556304 291796
rect 556264 6914 556292 291790
rect 557552 16574 557580 556407
rect 560312 16574 560340 557495
rect 565084 404388 565136 404394
rect 565084 404330 565136 404336
rect 562324 358828 562376 358834
rect 562324 358770 562376 358776
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 556172 6886 556292 6914
rect 555424 3664 555476 3670
rect 555424 3606 555476 3612
rect 554964 3052 555016 3058
rect 554964 2994 555016 3000
rect 554976 480 555004 2994
rect 556172 480 556200 6886
rect 557356 3800 557408 3806
rect 557356 3742 557408 3748
rect 557368 480 557396 3742
rect 558564 480 558592 16546
rect 559746 6352 559802 6361
rect 559746 6287 559802 6296
rect 559760 480 559788 6287
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 354 560432 16546
rect 562048 7608 562100 7614
rect 562048 7550 562100 7556
rect 562060 480 562088 7550
rect 562336 3534 562364 358770
rect 565096 333946 565124 404330
rect 565084 333940 565136 333946
rect 565084 333882 565136 333888
rect 565832 16574 565860 557534
rect 568580 316736 568632 316742
rect 568580 316678 568632 316684
rect 567844 272536 567896 272542
rect 567844 272478 567896 272484
rect 565832 16546 566872 16574
rect 565636 3664 565688 3670
rect 565636 3606 565688 3612
rect 563244 3596 563296 3602
rect 563244 3538 563296 3544
rect 562324 3528 562376 3534
rect 562324 3470 562376 3476
rect 563256 480 563284 3538
rect 564440 3460 564492 3466
rect 564440 3402 564492 3408
rect 564452 480 564480 3402
rect 565648 480 565676 3606
rect 566844 480 566872 16546
rect 567856 3330 567884 272478
rect 568592 16574 568620 316678
rect 569972 16574 570000 561682
rect 571984 556232 572036 556238
rect 571984 556174 572036 556180
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 568026 3496 568082 3505
rect 568026 3431 568082 3440
rect 567844 3324 567896 3330
rect 567844 3266 567896 3272
rect 568040 480 568068 3431
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 571996 3330 572024 556174
rect 572824 16574 572852 561886
rect 576124 561876 576176 561882
rect 576124 561818 576176 561824
rect 574100 551336 574152 551342
rect 574100 551278 574152 551284
rect 574112 16574 574140 551278
rect 572824 16546 573496 16574
rect 574112 16546 575152 16574
rect 571524 3324 571576 3330
rect 571524 3266 571576 3272
rect 571984 3324 572036 3330
rect 571984 3266 572036 3272
rect 572720 3324 572772 3330
rect 572720 3266 572772 3272
rect 571536 480 571564 3266
rect 572732 480 572760 3266
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576136 3398 576164 561818
rect 580356 555484 580408 555490
rect 580356 555426 580408 555432
rect 580264 554056 580316 554062
rect 580264 553998 580316 554004
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579618 471472 579674 471481
rect 579618 471407 579674 471416
rect 579632 470626 579660 471407
rect 579620 470620 579672 470626
rect 579620 470562 579672 470568
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 429894 580212 431559
rect 580172 429888 580224 429894
rect 580172 429830 580224 429836
rect 579710 418296 579766 418305
rect 579710 418231 579766 418240
rect 579724 418198 579752 418231
rect 579712 418192 579764 418198
rect 579712 418134 579764 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 578238 330440 578294 330449
rect 578238 330375 578294 330384
rect 578252 16574 578280 330375
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580276 219065 580304 553998
rect 580368 232393 580396 555426
rect 580446 524512 580502 524521
rect 580446 524447 580502 524456
rect 580460 338094 580488 524447
rect 580538 458144 580594 458153
rect 580538 458079 580594 458088
rect 580448 338088 580500 338094
rect 580448 338030 580500 338036
rect 580552 338026 580580 458079
rect 580630 351928 580686 351937
rect 580630 351863 580686 351872
rect 580540 338020 580592 338026
rect 580540 337962 580592 337968
rect 580644 337482 580672 351863
rect 580632 337476 580684 337482
rect 580632 337418 580684 337424
rect 580998 318064 581054 318073
rect 580998 317999 581054 318008
rect 580632 301504 580684 301510
rect 580632 301446 580684 301452
rect 580644 258913 580672 301446
rect 580630 258904 580686 258913
rect 580630 258839 580686 258848
rect 580446 258768 580502 258777
rect 580446 258703 580502 258712
rect 580354 232384 580410 232393
rect 580354 232319 580410 232328
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 579988 206984 580040 206990
rect 579988 206926 580040 206932
rect 580000 205737 580028 206926
rect 579986 205728 580042 205737
rect 579986 205663 580042 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579988 153196 580040 153202
rect 579988 153138 580040 153144
rect 580000 152697 580028 153138
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580264 138712 580316 138718
rect 580264 138654 580316 138660
rect 580276 126041 580304 138654
rect 580262 126032 580318 126041
rect 580262 125967 580318 125976
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580460 59673 580488 258703
rect 580446 59664 580502 59673
rect 580446 59599 580502 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 578252 16546 578648 16574
rect 576308 3528 576360 3534
rect 576308 3470 576360 3476
rect 576124 3392 576176 3398
rect 576124 3334 576176 3340
rect 576320 480 576348 3470
rect 577412 3392 577464 3398
rect 577412 3334 577464 3340
rect 577424 480 577452 3334
rect 578620 480 578648 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581012 480 581040 317999
rect 581090 279440 581146 279449
rect 581090 279375 581146 279384
rect 581104 16574 581132 279375
rect 581104 16546 581776 16574
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3146 619112 3202 619168
rect 3422 606056 3478 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3330 553832 3386 553888
rect 18 320728 74 320784
rect 3330 527856 3386 527912
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3238 501744 3294 501800
rect 3330 475668 3332 475688
rect 3332 475668 3384 475688
rect 3384 475668 3386 475688
rect 3330 475632 3386 475668
rect 3330 449520 3386 449576
rect 3146 423544 3202 423600
rect 3330 410488 3386 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 345344 3386 345400
rect 3146 254088 3202 254144
rect 3606 462576 3662 462632
rect 3514 371320 3570 371376
rect 3514 358400 3570 358456
rect 3514 319232 3570 319288
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 3514 267144 3570 267200
rect 3422 241032 3478 241088
rect 3330 214920 3386 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 2870 166232 2926 166288
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 5538 327664 5594 327720
rect 8298 553968 8354 554024
rect 11058 557096 11114 557152
rect 3422 6432 3478 6488
rect 19338 333240 19394 333296
rect 37278 558184 37334 558240
rect 22098 312432 22154 312488
rect 20626 3304 20682 3360
rect 32402 3440 32458 3496
rect 35898 322088 35954 322144
rect 45558 556960 45614 557016
rect 41418 313928 41474 313984
rect 39578 3576 39634 3632
rect 44270 316648 44326 316704
rect 56598 309712 56654 309768
rect 63498 333376 63554 333432
rect 60830 314064 60886 314120
rect 64878 251776 64934 251832
rect 71778 315288 71834 315344
rect 75918 320864 75974 320920
rect 93858 283464 93914 283520
rect 97998 311072 98054 311128
rect 93950 15816 94006 15872
rect 110418 323584 110474 323640
rect 118790 295976 118846 296032
rect 124218 333512 124274 333568
rect 135258 301416 135314 301472
rect 140778 557640 140834 557696
rect 138846 3848 138902 3904
rect 146298 335960 146354 336016
rect 154578 112376 154634 112432
rect 157338 334600 157394 334656
rect 171138 336096 171194 336152
rect 186318 336368 186374 336424
rect 182178 336232 182234 336288
rect 180798 308352 180854 308408
rect 179050 3984 179106 4040
rect 184938 11600 184994 11656
rect 212538 323720 212594 323776
rect 213826 6432 213882 6488
rect 220082 559000 220138 559056
rect 220450 338952 220506 339008
rect 223302 6568 223358 6624
rect 225694 559544 225750 559600
rect 224866 555872 224922 555928
rect 224406 6160 224462 6216
rect 224774 3712 224830 3768
rect 225694 338544 225750 338600
rect 226798 338680 226854 338736
rect 229834 554784 229890 554840
rect 228454 339224 228510 339280
rect 232042 555600 232098 555656
rect 232042 554240 232098 554296
rect 232042 552880 232098 552936
rect 232042 551520 232098 551576
rect 231674 548800 231730 548856
rect 231582 509360 231638 509416
rect 229926 338816 229982 338872
rect 231398 479440 231454 479496
rect 231306 476720 231362 476776
rect 231214 431840 231270 431896
rect 231122 389680 231178 389736
rect 230478 333104 230534 333160
rect 231490 448840 231546 448896
rect 232686 559680 232742 559736
rect 232594 559408 232650 559464
rect 232502 555192 232558 555248
rect 232042 546080 232098 546136
rect 232042 542000 232098 542056
rect 232042 539960 232098 540016
rect 232042 538600 232098 538656
rect 232042 537240 232098 537296
rect 232042 534520 232098 534576
rect 232318 533160 232374 533216
rect 232042 530440 232098 530496
rect 232042 529080 232098 529136
rect 232042 526360 232098 526416
rect 232042 525000 232098 525056
rect 232042 522280 232098 522336
rect 232042 520276 232044 520296
rect 232044 520276 232096 520296
rect 232096 520276 232098 520296
rect 232042 520240 232098 520276
rect 232042 518916 232044 518936
rect 232044 518916 232096 518936
rect 232096 518916 232098 518936
rect 232042 518880 232098 518916
rect 232042 516180 232098 516216
rect 232042 516160 232044 516180
rect 232044 516160 232096 516180
rect 232096 516160 232098 516180
rect 232042 510720 232098 510776
rect 231766 508000 231822 508056
rect 232042 506640 232098 506696
rect 232042 505280 232098 505336
rect 232042 502560 232098 502616
rect 232042 501200 232098 501256
rect 232042 496440 232098 496496
rect 232042 489640 232098 489696
rect 231858 486920 231914 486976
rect 232042 485560 232098 485616
rect 232042 482840 232098 482896
rect 232042 481480 232098 481536
rect 232042 478080 232098 478136
rect 232042 475360 232098 475416
rect 231858 474000 231914 474056
rect 232042 472640 232098 472696
rect 232042 471280 232098 471336
rect 232042 465840 232098 465896
rect 232042 464480 232098 464536
rect 232042 463120 232098 463176
rect 232042 461760 232098 461816
rect 232042 460400 232098 460456
rect 231950 458360 232006 458416
rect 232042 457000 232098 457056
rect 231950 455640 232006 455696
rect 232042 454280 232098 454336
rect 232042 452920 232098 452976
rect 232042 451560 232098 451616
rect 232318 444760 232374 444816
rect 232042 443400 232098 443456
rect 232042 442040 232098 442096
rect 232042 440680 232098 440736
rect 231950 434560 232006 434616
rect 232042 433236 232044 433256
rect 232044 433236 232096 433256
rect 232096 433236 232098 433256
rect 232042 433200 232098 433236
rect 231858 430480 231914 430536
rect 232042 429120 232098 429176
rect 232042 426436 232044 426456
rect 232044 426436 232096 426456
rect 232096 426436 232098 426456
rect 232042 426400 232098 426436
rect 232042 425076 232044 425096
rect 232044 425076 232096 425096
rect 232096 425076 232098 425096
rect 232042 425040 232098 425076
rect 232042 423700 232098 423736
rect 232042 423680 232044 423700
rect 232044 423680 232096 423700
rect 232096 423680 232098 423700
rect 232042 419600 232098 419656
rect 231950 416200 232006 416256
rect 232042 413480 232098 413536
rect 232042 410760 232098 410816
rect 232042 408040 232098 408096
rect 232410 403960 232466 404016
rect 232042 402600 232098 402656
rect 232042 399880 232098 399936
rect 232042 397840 232098 397896
rect 231950 396480 232006 396536
rect 232042 395120 232098 395176
rect 232410 393760 232466 393816
rect 232042 391040 232098 391096
rect 232042 385600 232098 385656
rect 232042 384240 232098 384296
rect 232042 378800 232098 378856
rect 232134 376760 232190 376816
rect 232042 375420 232098 375456
rect 232042 375400 232044 375420
rect 232044 375400 232096 375420
rect 232096 375400 232098 375420
rect 231858 374060 231914 374096
rect 231858 374040 231860 374060
rect 231860 374040 231912 374060
rect 231912 374040 231914 374060
rect 232042 372680 232098 372736
rect 232042 371320 232098 371376
rect 232042 368600 232098 368656
rect 231858 367240 231914 367296
rect 232042 363160 232098 363216
rect 232042 361800 232098 361856
rect 232042 357040 232098 357096
rect 232042 352960 232098 353016
rect 232042 351600 232098 351656
rect 232042 350240 232098 350296
rect 232042 348880 232098 348936
rect 232042 346160 232098 346216
rect 231950 344800 232006 344856
rect 232042 343440 232098 343496
rect 231950 342080 232006 342136
rect 232042 340720 232098 340776
rect 232042 339360 232098 339416
rect 232318 354320 232374 354376
rect 232226 339904 232282 339960
rect 230110 6296 230166 6352
rect 233054 556008 233110 556064
rect 232870 493720 232926 493776
rect 232870 450200 232926 450256
rect 232594 435920 232650 435976
rect 232502 364520 232558 364576
rect 232778 422320 232834 422376
rect 232686 382880 232742 382936
rect 232594 347520 232650 347576
rect 232502 339768 232558 339824
rect 233146 495080 233202 495136
rect 233054 412120 233110 412176
rect 233790 380160 233846 380216
rect 233606 359080 233662 359136
rect 233698 355680 233754 355736
rect 234066 555056 234122 555112
rect 234158 484200 234214 484256
rect 234250 468560 234306 468616
rect 234250 438640 234306 438696
rect 234066 420960 234122 421016
rect 233974 392400 234030 392456
rect 233882 360440 233938 360496
rect 234158 401240 234214 401296
rect 234434 555464 234490 555520
rect 234342 409400 234398 409456
rect 234342 405320 234398 405376
rect 234250 338136 234306 338192
rect 234526 547440 234582 547496
rect 234526 499160 234582 499216
rect 234434 358400 234490 358456
rect 234802 559136 234858 559192
rect 243404 556552 243460 556608
rect 251086 557504 251142 557560
rect 277858 557776 277914 557832
rect 282044 556824 282100 556880
rect 299432 556824 299488 556880
rect 304906 559272 304962 559328
rect 327078 557096 327134 557152
rect 330666 558048 330722 558104
rect 347962 560496 348018 560552
rect 346766 559816 346822 559872
rect 358358 559816 358414 559872
rect 365810 559680 365866 559736
rect 367006 558184 367062 558240
rect 375378 559544 375434 559600
rect 373170 556960 373226 557016
rect 384118 559408 384174 559464
rect 414938 560360 414994 560416
rect 409234 559000 409290 559056
rect 410522 557912 410578 557968
rect 417606 559136 417662 559192
rect 429198 557640 429254 557696
rect 440790 559544 440846 559600
rect 439502 559136 439558 559192
rect 444286 559408 444342 559464
rect 448426 559000 448482 559056
rect 450772 556688 450828 556744
rect 313600 556416 313656 556472
rect 319396 556416 319452 556472
rect 325836 556280 325892 556336
rect 235032 556008 235088 556064
rect 236320 555872 236376 555928
rect 264656 555872 264712 555928
rect 338072 555872 338128 555928
rect 352240 555872 352296 555928
rect 234710 417560 234766 417616
rect 234802 369960 234858 370016
rect 240506 338136 240562 338192
rect 267738 338136 267794 338192
rect 270774 338136 270830 338192
rect 379518 338136 379574 338192
rect 398930 338136 398986 338192
rect 412362 338136 412418 338192
rect 237378 337864 237434 337920
rect 238758 337592 238814 337648
rect 266358 327800 266414 327856
rect 302238 336504 302294 336560
rect 310242 6568 310298 6624
rect 316038 336640 316094 336696
rect 318798 337456 318854 337512
rect 327998 3848 328054 3904
rect 329194 3168 329250 3224
rect 337474 3984 337530 4040
rect 351642 3984 351698 4040
rect 356334 6432 356390 6488
rect 358818 337456 358874 337512
rect 363050 3440 363106 3496
rect 364430 3576 364486 3632
rect 367742 337320 367798 337376
rect 365810 6432 365866 6488
rect 381542 3304 381598 3360
rect 382370 316920 382426 316976
rect 390558 326304 390614 326360
rect 391846 3440 391902 3496
rect 441618 334056 441674 334112
rect 436742 3576 436798 3632
rect 437938 3168 437994 3224
rect 445758 304136 445814 304192
rect 450358 338136 450414 338192
rect 449898 337592 449954 337648
rect 447782 293120 447838 293176
rect 451646 513440 451702 513496
rect 451738 495080 451794 495136
rect 452934 559816 452990 559872
rect 452750 555056 452806 555112
rect 452658 491000 452714 491056
rect 451830 480120 451886 480176
rect 452106 474000 452162 474056
rect 452014 457680 452070 457736
rect 452658 468580 452714 468616
rect 452658 468560 452660 468580
rect 452660 468560 452712 468580
rect 452712 468560 452714 468580
rect 452658 459040 452714 459096
rect 452842 531800 452898 531856
rect 452750 430480 452806 430536
rect 452750 423680 452806 423736
rect 452842 409944 452898 410000
rect 452658 409400 452714 409456
rect 452658 401240 452714 401296
rect 452198 391040 452254 391096
rect 452842 388320 452898 388376
rect 452750 374720 452806 374776
rect 452658 355000 452714 355056
rect 453210 508000 453266 508056
rect 453210 482840 453266 482896
rect 453210 464480 453266 464536
rect 453026 451560 453082 451616
rect 453026 447500 453082 447536
rect 453026 447480 453028 447500
rect 453028 447480 453080 447500
rect 453080 447480 453082 447500
rect 453026 427760 453082 427816
rect 452934 344800 452990 344856
rect 453210 416900 453266 416936
rect 453210 416880 453212 416900
rect 453212 416880 453264 416900
rect 453264 416880 453266 416900
rect 453210 382900 453266 382936
rect 453210 382880 453212 382900
rect 453212 382880 453264 382900
rect 453264 382880 453266 382900
rect 453118 380160 453174 380216
rect 453394 550160 453450 550216
rect 453946 554240 454002 554296
rect 453946 547440 454002 547496
rect 453946 546080 454002 546136
rect 453578 544720 453634 544776
rect 453946 543360 454002 543416
rect 453762 542000 453818 542056
rect 453762 537920 453818 537976
rect 453946 535880 454002 535936
rect 453946 533160 454002 533216
rect 453578 530440 453634 530496
rect 453946 527720 454002 527776
rect 453670 525000 453726 525056
rect 453946 522280 454002 522336
rect 453946 520940 454002 520976
rect 453946 520920 453948 520940
rect 453948 520920 454000 520940
rect 454000 520920 454002 520940
rect 453946 519560 454002 519616
rect 453946 514820 454002 514856
rect 453946 514800 453948 514820
rect 453948 514800 454000 514820
rect 454000 514800 454002 514820
rect 453762 512080 453818 512136
rect 453762 509360 453818 509416
rect 453946 503920 454002 503976
rect 453578 502560 453634 502616
rect 453946 499840 454002 499896
rect 453946 498500 454002 498536
rect 453946 498480 453948 498500
rect 453948 498480 454000 498500
rect 454000 498480 454002 498500
rect 453946 492360 454002 492416
rect 453762 489640 453818 489696
rect 453946 488280 454002 488336
rect 453762 486920 453818 486976
rect 453946 485560 454002 485616
rect 453762 481480 453818 481536
rect 453762 478760 453818 478816
rect 453854 477400 453910 477456
rect 453946 476040 454002 476096
rect 453946 472640 454002 472696
rect 453762 471300 453818 471336
rect 453762 471280 453764 471300
rect 453764 471280 453816 471300
rect 453816 471280 453818 471300
rect 453946 469920 454002 469976
rect 453578 467200 453634 467256
rect 453946 463120 454002 463176
rect 453946 460400 454002 460456
rect 453670 456320 453726 456376
rect 453946 454300 454002 454336
rect 453946 454280 453948 454300
rect 453948 454280 454000 454300
rect 454000 454280 454002 454300
rect 453946 452920 454002 452976
rect 453578 450220 453634 450256
rect 453578 450200 453580 450220
rect 453580 450200 453632 450220
rect 453632 450200 453634 450220
rect 453946 444780 454002 444816
rect 453946 444760 453948 444780
rect 453948 444760 454000 444780
rect 454000 444760 454002 444780
rect 453946 440680 454002 440736
rect 453854 439320 453910 439376
rect 453946 437960 454002 438016
rect 453946 436600 454002 436656
rect 453670 435240 453726 435296
rect 453946 431840 454002 431896
rect 453946 429120 454002 429176
rect 453946 426436 453948 426456
rect 453948 426436 454000 426456
rect 454000 426436 454002 426456
rect 453946 426400 454002 426436
rect 453946 425076 453948 425096
rect 453948 425076 454000 425096
rect 454000 425076 454002 425096
rect 453946 425040 454002 425076
rect 453946 420980 454002 421016
rect 453946 420960 453948 420980
rect 453948 420960 454000 420980
rect 454000 420960 454002 420980
rect 453670 418260 453726 418296
rect 453670 418240 453672 418260
rect 453672 418240 453724 418260
rect 453724 418240 453726 418260
rect 453946 413480 454002 413536
rect 453762 408040 453818 408096
rect 453946 406680 454002 406736
rect 453762 405320 453818 405376
rect 453946 402600 454002 402656
rect 453762 399880 453818 399936
rect 453762 395800 453818 395856
rect 453762 394440 453818 394496
rect 453946 392400 454002 392456
rect 453946 389680 454002 389736
rect 453946 386960 454002 387016
rect 453946 385636 453948 385656
rect 453948 385636 454000 385656
rect 454000 385636 454002 385656
rect 453946 385600 454002 385636
rect 453946 384240 454002 384296
rect 453762 378820 453818 378856
rect 453762 378800 453764 378820
rect 453764 378800 453816 378820
rect 453816 378800 453818 378820
rect 453762 376080 453818 376136
rect 453946 372700 454002 372736
rect 453946 372680 453948 372700
rect 453948 372680 454000 372700
rect 454000 372680 454002 372700
rect 453762 371320 453818 371376
rect 453762 369960 453818 370016
rect 453762 368600 453818 368656
rect 453946 367260 454002 367296
rect 453946 367240 453948 367260
rect 453948 367240 454000 367260
rect 454000 367240 454002 367260
rect 453946 365880 454002 365936
rect 453762 364520 453818 364576
rect 453762 363160 453818 363216
rect 453578 356360 453634 356416
rect 453486 353640 453542 353696
rect 453210 346160 453266 346216
rect 453670 350240 453726 350296
rect 453578 338272 453634 338328
rect 453946 361800 454002 361856
rect 453946 359080 454002 359136
rect 453946 357720 454002 357776
rect 453946 348880 454002 348936
rect 454130 526360 454186 526416
rect 453946 347556 453948 347576
rect 453948 347556 454000 347576
rect 454000 347556 454002 347576
rect 453946 347520 454002 347556
rect 453946 343440 454002 343496
rect 453946 342100 454002 342136
rect 453946 342080 453948 342100
rect 453948 342080 454000 342100
rect 454000 342080 454002 342100
rect 454038 341400 454094 341456
rect 454222 465840 454278 465896
rect 456798 300056 456854 300112
rect 456890 261432 456946 261488
rect 457074 338816 457130 338872
rect 457534 339224 457590 339280
rect 458362 339632 458418 339688
rect 458822 338544 458878 338600
rect 458914 333376 458970 333432
rect 460110 335960 460166 336016
rect 460386 338680 460442 338736
rect 463790 559272 463846 559328
rect 461674 338952 461730 339008
rect 463974 559136 464030 559192
rect 463974 337456 464030 337512
rect 463790 3168 463846 3224
rect 465262 559408 465318 559464
rect 465446 336368 465502 336424
rect 465538 333240 465594 333296
rect 465262 36488 465318 36544
rect 474002 559544 474058 559600
rect 465906 3576 465962 3632
rect 476118 37848 476174 37904
rect 505098 331744 505154 331800
rect 507858 329160 507914 329216
rect 517518 329024 517574 329080
rect 523130 316784 523186 316840
rect 521658 170312 521714 170368
rect 530122 3712 530178 3768
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580354 577632 580410 577688
rect 579802 564304 579858 564360
rect 560298 557504 560354 557560
rect 557538 556416 557594 556472
rect 550638 556280 550694 556336
rect 552018 318144 552074 318200
rect 553766 6160 553822 6216
rect 559746 6296 559802 6352
rect 568026 3440 568082 3496
rect 580170 537784 580226 537840
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579618 471416 579674 471472
rect 580170 431568 580226 431624
rect 579710 418240 579766 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 578238 330384 578294 330440
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580446 524456 580502 524512
rect 580538 458088 580594 458144
rect 580630 351872 580686 351928
rect 580998 318008 581054 318064
rect 580630 258848 580686 258904
rect 580446 258712 580502 258768
rect 580354 232328 580410 232384
rect 580262 219000 580318 219056
rect 579986 205672 580042 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 579986 152632 580042 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580262 125976 580318 126032
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580446 59608 580502 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
rect 581090 279384 581146 279440
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 460974 632090 460980 632092
rect -960 632030 460980 632090
rect -960 631940 480 632030
rect 460974 632028 460980 632030
rect 461044 632028 461050 632092
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580349 577690 580415 577693
rect 583520 577690 584960 577780
rect 580349 577688 584960 577690
rect 580349 577632 580354 577688
rect 580410 577632 584960 577688
rect 580349 577630 584960 577632
rect 580349 577627 580415 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect 225638 560492 225644 560556
rect 225708 560554 225714 560556
rect 347957 560554 348023 560557
rect 225708 560552 348023 560554
rect 225708 560496 347962 560552
rect 348018 560496 348023 560552
rect 225708 560494 348023 560496
rect 225708 560492 225714 560494
rect 347957 560491 348023 560494
rect 227110 560356 227116 560420
rect 227180 560418 227186 560420
rect 414933 560418 414999 560421
rect 227180 560416 414999 560418
rect 227180 560360 414938 560416
rect 414994 560360 414999 560416
rect 227180 560358 414999 560360
rect 227180 560356 227186 560358
rect 414933 560355 414999 560358
rect 226190 559812 226196 559876
rect 226260 559874 226266 559876
rect 346761 559874 346827 559877
rect 226260 559872 346827 559874
rect 226260 559816 346766 559872
rect 346822 559816 346827 559872
rect 226260 559814 346827 559816
rect 226260 559812 226266 559814
rect 346761 559811 346827 559814
rect 358353 559874 358419 559877
rect 452929 559874 452995 559877
rect 358353 559872 452995 559874
rect 358353 559816 358358 559872
rect 358414 559816 452934 559872
rect 452990 559816 452995 559872
rect 358353 559814 452995 559816
rect 358353 559811 358419 559814
rect 452929 559811 452995 559814
rect 232681 559738 232747 559741
rect 365805 559738 365871 559741
rect 232681 559736 365871 559738
rect 232681 559680 232686 559736
rect 232742 559680 365810 559736
rect 365866 559680 365871 559736
rect 232681 559678 365871 559680
rect 232681 559675 232747 559678
rect 365805 559675 365871 559678
rect 225689 559602 225755 559605
rect 375373 559602 375439 559605
rect 225689 559600 375439 559602
rect 225689 559544 225694 559600
rect 225750 559544 375378 559600
rect 375434 559544 375439 559600
rect 225689 559542 375439 559544
rect 225689 559539 225755 559542
rect 375373 559539 375439 559542
rect 440785 559602 440851 559605
rect 473997 559602 474063 559605
rect 440785 559600 474063 559602
rect 440785 559544 440790 559600
rect 440846 559544 474002 559600
rect 474058 559544 474063 559600
rect 440785 559542 474063 559544
rect 440785 559539 440851 559542
rect 473997 559539 474063 559542
rect 232589 559466 232655 559469
rect 384113 559466 384179 559469
rect 232589 559464 384179 559466
rect 232589 559408 232594 559464
rect 232650 559408 384118 559464
rect 384174 559408 384179 559464
rect 232589 559406 384179 559408
rect 232589 559403 232655 559406
rect 384113 559403 384179 559406
rect 444281 559466 444347 559469
rect 465257 559466 465323 559469
rect 444281 559464 465323 559466
rect 444281 559408 444286 559464
rect 444342 559408 465262 559464
rect 465318 559408 465323 559464
rect 444281 559406 465323 559408
rect 444281 559403 444347 559406
rect 465257 559403 465323 559406
rect 304901 559330 304967 559333
rect 463785 559330 463851 559333
rect 304901 559328 463851 559330
rect 304901 559272 304906 559328
rect 304962 559272 463790 559328
rect 463846 559272 463851 559328
rect 304901 559270 463851 559272
rect 304901 559267 304967 559270
rect 463785 559267 463851 559270
rect 234797 559194 234863 559197
rect 417601 559194 417667 559197
rect 234797 559192 417667 559194
rect 234797 559136 234802 559192
rect 234858 559136 417606 559192
rect 417662 559136 417667 559192
rect 234797 559134 417667 559136
rect 234797 559131 234863 559134
rect 417601 559131 417667 559134
rect 439497 559194 439563 559197
rect 463969 559194 464035 559197
rect 439497 559192 464035 559194
rect 439497 559136 439502 559192
rect 439558 559136 463974 559192
rect 464030 559136 464035 559192
rect 439497 559134 464035 559136
rect 439497 559131 439563 559134
rect 463969 559131 464035 559134
rect 220077 559058 220143 559061
rect 409229 559058 409295 559061
rect 220077 559056 409295 559058
rect 220077 559000 220082 559056
rect 220138 559000 409234 559056
rect 409290 559000 409295 559056
rect 220077 558998 409295 559000
rect 220077 558995 220143 558998
rect 409229 558995 409295 558998
rect 448421 559058 448487 559061
rect 461158 559058 461164 559060
rect 448421 559056 461164 559058
rect 448421 559000 448426 559056
rect 448482 559000 461164 559056
rect 448421 558998 461164 559000
rect 448421 558995 448487 558998
rect 461158 558996 461164 558998
rect 461228 558996 461234 559060
rect 37273 558242 37339 558245
rect 367001 558242 367067 558245
rect 37273 558240 367067 558242
rect 37273 558184 37278 558240
rect 37334 558184 367006 558240
rect 367062 558184 367067 558240
rect 37273 558182 367067 558184
rect 37273 558179 37339 558182
rect 367001 558179 367067 558182
rect 229686 558044 229692 558108
rect 229756 558106 229762 558108
rect 330661 558106 330727 558109
rect 229756 558104 330727 558106
rect 229756 558048 330666 558104
rect 330722 558048 330727 558104
rect 229756 558046 330727 558048
rect 229756 558044 229762 558046
rect 330661 558043 330727 558046
rect 228214 557908 228220 557972
rect 228284 557970 228290 557972
rect 410517 557970 410583 557973
rect 228284 557968 410583 557970
rect 228284 557912 410522 557968
rect 410578 557912 410583 557968
rect 228284 557910 410583 557912
rect 228284 557908 228290 557910
rect 410517 557907 410583 557910
rect 277853 557834 277919 557837
rect 460054 557834 460060 557836
rect 277853 557832 460060 557834
rect 277853 557776 277858 557832
rect 277914 557776 460060 557832
rect 277853 557774 460060 557776
rect 277853 557771 277919 557774
rect 460054 557772 460060 557774
rect 460124 557772 460130 557836
rect 140773 557698 140839 557701
rect 429193 557698 429259 557701
rect 140773 557696 429259 557698
rect 140773 557640 140778 557696
rect 140834 557640 429198 557696
rect 429254 557640 429259 557696
rect 140773 557638 429259 557640
rect 140773 557635 140839 557638
rect 429193 557635 429259 557638
rect 251081 557562 251147 557565
rect 560293 557562 560359 557565
rect 251081 557560 560359 557562
rect 251081 557504 251086 557560
rect 251142 557504 560298 557560
rect 560354 557504 560359 557560
rect 251081 557502 560359 557504
rect 251081 557499 251147 557502
rect 560293 557499 560359 557502
rect 11053 557154 11119 557157
rect 327073 557154 327139 557157
rect 11053 557152 327139 557154
rect 11053 557096 11058 557152
rect 11114 557096 327078 557152
rect 327134 557096 327139 557152
rect 11053 557094 327139 557096
rect 11053 557091 11119 557094
rect 327073 557091 327139 557094
rect 45553 557018 45619 557021
rect 373165 557018 373231 557021
rect 45553 557016 373231 557018
rect 45553 556960 45558 557016
rect 45614 556960 373170 557016
rect 373226 556960 373231 557016
rect 45553 556958 373231 556960
rect 45553 556955 45619 556958
rect 373165 556955 373231 556958
rect 228950 556820 228956 556884
rect 229020 556882 229026 556884
rect 282039 556882 282105 556885
rect 229020 556880 282105 556882
rect 229020 556824 282044 556880
rect 282100 556824 282105 556880
rect 229020 556822 282105 556824
rect 229020 556820 229026 556822
rect 282039 556819 282105 556822
rect 299427 556882 299493 556885
rect 451038 556882 451044 556884
rect 299427 556880 451044 556882
rect 299427 556824 299432 556880
rect 299488 556824 451044 556880
rect 299427 556822 451044 556824
rect 299427 556819 299493 556822
rect 451038 556820 451044 556822
rect 451108 556820 451114 556884
rect 235758 556684 235764 556748
rect 235828 556746 235834 556748
rect 450767 556746 450833 556749
rect 235828 556744 450833 556746
rect 235828 556688 450772 556744
rect 450828 556688 450833 556744
rect 235828 556686 450833 556688
rect 235828 556684 235834 556686
rect 450767 556683 450833 556686
rect 243399 556610 243465 556613
rect 460238 556610 460244 556612
rect 243399 556608 460244 556610
rect 243399 556552 243404 556608
rect 243460 556552 460244 556608
rect 243399 556550 460244 556552
rect 243399 556547 243465 556550
rect 460238 556548 460244 556550
rect 460308 556548 460314 556612
rect 225454 556412 225460 556476
rect 225524 556474 225530 556476
rect 313595 556474 313661 556477
rect 225524 556472 313661 556474
rect 225524 556416 313600 556472
rect 313656 556416 313661 556472
rect 225524 556414 313661 556416
rect 225524 556412 225530 556414
rect 313595 556411 313661 556414
rect 319391 556474 319457 556477
rect 557533 556474 557599 556477
rect 319391 556472 557599 556474
rect 319391 556416 319396 556472
rect 319452 556416 557538 556472
rect 557594 556416 557599 556472
rect 319391 556414 557599 556416
rect 319391 556411 319457 556414
rect 557533 556411 557599 556414
rect 325831 556338 325897 556341
rect 550633 556338 550699 556341
rect 325831 556336 550699 556338
rect 325831 556280 325836 556336
rect 325892 556280 550638 556336
rect 550694 556280 550699 556336
rect 325831 556278 550699 556280
rect 325831 556275 325897 556278
rect 550633 556275 550699 556278
rect 233049 556066 233115 556069
rect 235027 556066 235093 556069
rect 233049 556064 235093 556066
rect 233049 556008 233054 556064
rect 233110 556008 235032 556064
rect 235088 556008 235093 556064
rect 233049 556006 235093 556008
rect 233049 556003 233115 556006
rect 235027 556003 235093 556006
rect 224861 555930 224927 555933
rect 236315 555930 236381 555933
rect 264651 555932 264717 555933
rect 264646 555930 264652 555932
rect 224861 555928 236381 555930
rect 224861 555872 224866 555928
rect 224922 555872 236320 555928
rect 236376 555872 236381 555928
rect 224861 555870 236381 555872
rect 264560 555870 264652 555930
rect 224861 555867 224927 555870
rect 236315 555867 236381 555870
rect 264646 555868 264652 555870
rect 264716 555868 264722 555932
rect 338067 555930 338133 555933
rect 352235 555932 352301 555933
rect 352230 555930 352236 555932
rect 315990 555928 338133 555930
rect 315990 555872 338072 555928
rect 338128 555872 338133 555928
rect 315990 555870 338133 555872
rect 352144 555870 352236 555930
rect 264651 555867 264717 555868
rect 232037 555658 232103 555661
rect 232037 555656 235060 555658
rect 232037 555600 232042 555656
rect 232098 555600 235060 555656
rect 232037 555598 235060 555600
rect 232037 555595 232103 555598
rect 234429 555522 234495 555525
rect 315990 555522 316050 555870
rect 338067 555867 338133 555870
rect 352230 555868 352236 555870
rect 352300 555868 352306 555932
rect 352235 555867 352301 555868
rect 234429 555520 316050 555522
rect 234429 555464 234434 555520
rect 234490 555464 316050 555520
rect 234429 555462 316050 555464
rect 234429 555459 234495 555462
rect 232497 555250 232563 555253
rect 264646 555250 264652 555252
rect 232497 555248 264652 555250
rect 232497 555192 232502 555248
rect 232558 555192 264652 555248
rect 232497 555190 264652 555192
rect 232497 555187 232563 555190
rect 264646 555188 264652 555190
rect 264716 555188 264722 555252
rect 234061 555114 234127 555117
rect 452745 555114 452811 555117
rect 234061 555112 452811 555114
rect 234061 555056 234066 555112
rect 234122 555056 452750 555112
rect 452806 555056 452811 555112
rect 234061 555054 452811 555056
rect 234061 555051 234127 555054
rect 452745 555051 452811 555054
rect 229829 554842 229895 554845
rect 352230 554842 352236 554844
rect 229829 554840 352236 554842
rect 229829 554784 229834 554840
rect 229890 554784 352236 554840
rect 229829 554782 352236 554784
rect 229829 554779 229895 554782
rect 352230 554780 352236 554782
rect 352300 554780 352306 554844
rect 235758 554570 235764 554572
rect 219390 554510 235764 554570
rect 8293 554026 8359 554029
rect 219390 554026 219450 554510
rect 235758 554508 235764 554510
rect 235828 554508 235834 554572
rect 232037 554298 232103 554301
rect 453941 554298 454007 554301
rect 232037 554296 235060 554298
rect 232037 554240 232042 554296
rect 232098 554240 235060 554296
rect 232037 554238 235060 554240
rect 451444 554296 454007 554298
rect 451444 554240 453946 554296
rect 454002 554240 454007 554296
rect 451444 554238 454007 554240
rect 232037 554235 232103 554238
rect 453941 554235 454007 554238
rect 8293 554024 219450 554026
rect -960 553890 480 553980
rect 8293 553968 8298 554024
rect 8354 553968 219450 554024
rect 8293 553966 219450 553968
rect 8293 553963 8359 553966
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 232037 552938 232103 552941
rect 458398 552938 458404 552940
rect 232037 552936 235060 552938
rect 232037 552880 232042 552936
rect 232098 552880 235060 552936
rect 232037 552878 235060 552880
rect 451444 552878 458404 552938
rect 232037 552875 232103 552878
rect 458398 552876 458404 552878
rect 458468 552876 458474 552940
rect 232037 551578 232103 551581
rect 455638 551578 455644 551580
rect 232037 551576 235060 551578
rect 232037 551520 232042 551576
rect 232098 551520 235060 551576
rect 232037 551518 235060 551520
rect 451444 551518 455644 551578
rect 232037 551515 232103 551518
rect 455638 551516 455644 551518
rect 455708 551516 455714 551580
rect 583520 551020 584960 551260
rect 231158 550156 231164 550220
rect 231228 550218 231234 550220
rect 453389 550218 453455 550221
rect 231228 550158 235060 550218
rect 451444 550216 453455 550218
rect 451444 550160 453394 550216
rect 453450 550160 453455 550216
rect 451444 550158 453455 550160
rect 231228 550156 231234 550158
rect 453389 550155 453455 550158
rect 231669 548858 231735 548861
rect 458582 548858 458588 548860
rect 231669 548856 235060 548858
rect 231669 548800 231674 548856
rect 231730 548800 235060 548856
rect 231669 548798 235060 548800
rect 451444 548798 458588 548858
rect 231669 548795 231735 548798
rect 458582 548796 458588 548798
rect 458652 548796 458658 548860
rect 234521 547498 234587 547501
rect 453941 547498 454007 547501
rect 234521 547496 235060 547498
rect 234521 547440 234526 547496
rect 234582 547440 235060 547496
rect 234521 547438 235060 547440
rect 451444 547496 454007 547498
rect 451444 547440 453946 547496
rect 454002 547440 454007 547496
rect 451444 547438 454007 547440
rect 234521 547435 234587 547438
rect 453941 547435 454007 547438
rect 232037 546138 232103 546141
rect 453941 546138 454007 546141
rect 232037 546136 235060 546138
rect 232037 546080 232042 546136
rect 232098 546080 235060 546136
rect 232037 546078 235060 546080
rect 451444 546136 454007 546138
rect 451444 546080 453946 546136
rect 454002 546080 454007 546136
rect 451444 546078 454007 546080
rect 232037 546075 232103 546078
rect 453941 546075 454007 546078
rect 453573 544778 453639 544781
rect 451444 544776 453639 544778
rect 451444 544720 453578 544776
rect 453634 544720 453639 544776
rect 451444 544718 453639 544720
rect 453573 544715 453639 544718
rect 453941 543418 454007 543421
rect 451444 543416 454007 543418
rect 227294 542404 227300 542468
rect 227364 542466 227370 542468
rect 235030 542466 235090 543388
rect 451444 543360 453946 543416
rect 454002 543360 454007 543416
rect 451444 543358 454007 543360
rect 453941 543355 454007 543358
rect 227364 542406 235090 542466
rect 227364 542404 227370 542406
rect 232037 542058 232103 542061
rect 453757 542058 453823 542061
rect 232037 542056 235060 542058
rect 232037 542000 232042 542056
rect 232098 542000 235060 542056
rect 232037 541998 235060 542000
rect 451444 542056 453823 542058
rect 451444 542000 453762 542056
rect 453818 542000 453823 542056
rect 451444 541998 453823 542000
rect 232037 541995 232103 541998
rect 453757 541995 453823 541998
rect -960 540684 480 540924
rect 232037 540018 232103 540021
rect 232037 540016 235060 540018
rect 232037 539960 232042 540016
rect 232098 539960 235060 540016
rect 232037 539958 235060 539960
rect 232037 539955 232103 539958
rect 452878 539338 452884 539340
rect 451444 539278 452884 539338
rect 452878 539276 452884 539278
rect 452948 539276 452954 539340
rect 232037 538658 232103 538661
rect 232037 538656 235060 538658
rect 232037 538600 232042 538656
rect 232098 538600 235060 538656
rect 232037 538598 235060 538600
rect 232037 538595 232103 538598
rect 453757 537978 453823 537981
rect 451444 537976 453823 537978
rect 451444 537920 453762 537976
rect 453818 537920 453823 537976
rect 451444 537918 453823 537920
rect 453757 537915 453823 537918
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 232037 537298 232103 537301
rect 232037 537296 235060 537298
rect 232037 537240 232042 537296
rect 232098 537240 235060 537296
rect 232037 537238 235060 537240
rect 232037 537235 232103 537238
rect 231342 535876 231348 535940
rect 231412 535938 231418 535940
rect 453941 535938 454007 535941
rect 231412 535878 235060 535938
rect 451444 535936 454007 535938
rect 451444 535880 453946 535936
rect 454002 535880 454007 535936
rect 451444 535878 454007 535880
rect 231412 535876 231418 535878
rect 453941 535875 454007 535878
rect 232037 534578 232103 534581
rect 232037 534576 235060 534578
rect 232037 534520 232042 534576
rect 232098 534520 235060 534576
rect 232037 534518 235060 534520
rect 232037 534515 232103 534518
rect 232313 533218 232379 533221
rect 453941 533218 454007 533221
rect 232313 533216 235060 533218
rect 232313 533160 232318 533216
rect 232374 533160 235060 533216
rect 232313 533158 235060 533160
rect 451444 533216 454007 533218
rect 451444 533160 453946 533216
rect 454002 533160 454007 533216
rect 451444 533158 454007 533160
rect 232313 533155 232379 533158
rect 453941 533155 454007 533158
rect 452837 531858 452903 531861
rect 451444 531856 452903 531858
rect 227478 531388 227484 531452
rect 227548 531450 227554 531452
rect 235030 531450 235090 531828
rect 451444 531800 452842 531856
rect 452898 531800 452903 531856
rect 451444 531798 452903 531800
rect 452837 531795 452903 531798
rect 227548 531390 235090 531450
rect 227548 531388 227554 531390
rect 232037 530498 232103 530501
rect 453573 530498 453639 530501
rect 232037 530496 235060 530498
rect 232037 530440 232042 530496
rect 232098 530440 235060 530496
rect 232037 530438 235060 530440
rect 451444 530496 453639 530498
rect 451444 530440 453578 530496
rect 453634 530440 453639 530496
rect 451444 530438 453639 530440
rect 232037 530435 232103 530438
rect 453573 530435 453639 530438
rect 232037 529138 232103 529141
rect 458214 529138 458220 529140
rect 232037 529136 235060 529138
rect 232037 529080 232042 529136
rect 232098 529080 235060 529136
rect 232037 529078 235060 529080
rect 451444 529078 458220 529138
rect 232037 529075 232103 529078
rect 458214 529076 458220 529078
rect 458284 529076 458290 529140
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 230238 527716 230244 527780
rect 230308 527778 230314 527780
rect 453941 527778 454007 527781
rect 230308 527718 235060 527778
rect 451444 527776 454007 527778
rect 451444 527720 453946 527776
rect 454002 527720 454007 527776
rect 451444 527718 454007 527720
rect 230308 527716 230314 527718
rect 453941 527715 454007 527718
rect 232037 526418 232103 526421
rect 454125 526418 454191 526421
rect 232037 526416 235060 526418
rect 232037 526360 232042 526416
rect 232098 526360 235060 526416
rect 232037 526358 235060 526360
rect 451444 526416 454191 526418
rect 451444 526360 454130 526416
rect 454186 526360 454191 526416
rect 451444 526358 454191 526360
rect 232037 526355 232103 526358
rect 454125 526355 454191 526358
rect 232037 525058 232103 525061
rect 453665 525058 453731 525061
rect 232037 525056 235060 525058
rect 232037 525000 232042 525056
rect 232098 525000 235060 525056
rect 232037 524998 235060 525000
rect 451444 525056 453731 525058
rect 451444 525000 453670 525056
rect 453726 525000 453731 525056
rect 451444 524998 453731 525000
rect 232037 524995 232103 524998
rect 453665 524995 453731 524998
rect 580441 524514 580507 524517
rect 583520 524514 584960 524604
rect 580441 524512 584960 524514
rect 580441 524456 580446 524512
rect 580502 524456 584960 524512
rect 580441 524454 584960 524456
rect 580441 524451 580507 524454
rect 583520 524364 584960 524454
rect 233366 523636 233372 523700
rect 233436 523698 233442 523700
rect 456742 523698 456748 523700
rect 233436 523638 235060 523698
rect 451444 523638 456748 523698
rect 233436 523636 233442 523638
rect 456742 523636 456748 523638
rect 456812 523636 456818 523700
rect 232037 522338 232103 522341
rect 453941 522338 454007 522341
rect 232037 522336 235060 522338
rect 232037 522280 232042 522336
rect 232098 522280 235060 522336
rect 232037 522278 235060 522280
rect 451444 522336 454007 522338
rect 451444 522280 453946 522336
rect 454002 522280 454007 522336
rect 451444 522278 454007 522280
rect 232037 522275 232103 522278
rect 453941 522275 454007 522278
rect 453941 520978 454007 520981
rect 451444 520976 454007 520978
rect 451444 520920 453946 520976
rect 454002 520920 454007 520976
rect 451444 520918 454007 520920
rect 453941 520915 454007 520918
rect 232037 520298 232103 520301
rect 232037 520296 235060 520298
rect 232037 520240 232042 520296
rect 232098 520240 235060 520296
rect 232037 520238 235060 520240
rect 232037 520235 232103 520238
rect 453941 519618 454007 519621
rect 451444 519616 454007 519618
rect 451444 519560 453946 519616
rect 454002 519560 454007 519616
rect 451444 519558 454007 519560
rect 453941 519555 454007 519558
rect 232037 518938 232103 518941
rect 232037 518936 235060 518938
rect 232037 518880 232042 518936
rect 232098 518880 235060 518936
rect 232037 518878 235060 518880
rect 232037 518875 232103 518878
rect 228766 517516 228772 517580
rect 228836 517578 228842 517580
rect 228836 517518 235060 517578
rect 228836 517516 228842 517518
rect 232037 516218 232103 516221
rect 232037 516216 235060 516218
rect 232037 516160 232042 516216
rect 232098 516160 235060 516216
rect 232037 516158 235060 516160
rect 232037 516155 232103 516158
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect 453941 514858 454007 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect 451444 514856 454007 514858
rect 451444 514800 453946 514856
rect 454002 514800 454007 514856
rect 451444 514798 454007 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 453941 514795 454007 514798
rect 230054 513436 230060 513500
rect 230124 513498 230130 513500
rect 451641 513498 451707 513501
rect 230124 513438 235060 513498
rect 451444 513496 451707 513498
rect 451444 513440 451646 513496
rect 451702 513440 451707 513496
rect 451444 513438 451707 513440
rect 230124 513436 230130 513438
rect 451641 513435 451707 513438
rect 231710 512076 231716 512140
rect 231780 512138 231786 512140
rect 453757 512138 453823 512141
rect 231780 512078 235060 512138
rect 451444 512136 453823 512138
rect 451444 512080 453762 512136
rect 453818 512080 453823 512136
rect 451444 512078 453823 512080
rect 231780 512076 231786 512078
rect 453757 512075 453823 512078
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 232037 510778 232103 510781
rect 232037 510776 235060 510778
rect 232037 510720 232042 510776
rect 232098 510720 235060 510776
rect 232037 510718 235060 510720
rect 232037 510715 232103 510718
rect 451414 510642 451474 510748
rect 463734 510642 463740 510644
rect 451414 510582 463740 510642
rect 463734 510580 463740 510582
rect 463804 510580 463810 510644
rect 231577 509418 231643 509421
rect 453757 509418 453823 509421
rect 231577 509416 235060 509418
rect 231577 509360 231582 509416
rect 231638 509360 235060 509416
rect 231577 509358 235060 509360
rect 451444 509416 453823 509418
rect 451444 509360 453762 509416
rect 453818 509360 453823 509416
rect 451444 509358 453823 509360
rect 231577 509355 231643 509358
rect 453757 509355 453823 509358
rect 231761 508058 231827 508061
rect 453205 508058 453271 508061
rect 231761 508056 235060 508058
rect 231761 508000 231766 508056
rect 231822 508000 235060 508056
rect 231761 507998 235060 508000
rect 451444 508056 453271 508058
rect 451444 508000 453210 508056
rect 453266 508000 453271 508056
rect 451444 507998 453271 508000
rect 231761 507995 231827 507998
rect 453205 507995 453271 507998
rect 232037 506698 232103 506701
rect 232037 506696 235060 506698
rect 232037 506640 232042 506696
rect 232098 506640 235060 506696
rect 232037 506638 235060 506640
rect 232037 506635 232103 506638
rect 451414 506562 451474 506668
rect 461342 506562 461348 506564
rect 451414 506502 461348 506562
rect 461342 506500 461348 506502
rect 461412 506500 461418 506564
rect 232037 505338 232103 505341
rect 456926 505338 456932 505340
rect 232037 505336 235060 505338
rect 232037 505280 232042 505336
rect 232098 505280 235060 505336
rect 232037 505278 235060 505280
rect 451444 505278 456932 505338
rect 232037 505275 232103 505278
rect 456926 505276 456932 505278
rect 456996 505276 457002 505340
rect 233734 503916 233740 503980
rect 233804 503978 233810 503980
rect 453941 503978 454007 503981
rect 233804 503918 235060 503978
rect 451444 503976 454007 503978
rect 451444 503920 453946 503976
rect 454002 503920 454007 503976
rect 451444 503918 454007 503920
rect 233804 503916 233810 503918
rect 453941 503915 454007 503918
rect 232037 502618 232103 502621
rect 453573 502618 453639 502621
rect 232037 502616 235060 502618
rect 232037 502560 232042 502616
rect 232098 502560 235060 502616
rect 232037 502558 235060 502560
rect 451444 502616 453639 502618
rect 451444 502560 453578 502616
rect 453634 502560 453639 502616
rect 451444 502558 453639 502560
rect 232037 502555 232103 502558
rect 453573 502555 453639 502558
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 232037 501258 232103 501261
rect 458766 501258 458772 501260
rect 232037 501256 235060 501258
rect 232037 501200 232042 501256
rect 232098 501200 235060 501256
rect 232037 501198 235060 501200
rect 451444 501198 458772 501258
rect 232037 501195 232103 501198
rect 458766 501196 458772 501198
rect 458836 501196 458842 501260
rect 453941 499898 454007 499901
rect 451444 499896 454007 499898
rect 451444 499840 453946 499896
rect 454002 499840 454007 499896
rect 451444 499838 454007 499840
rect 453941 499835 454007 499838
rect 234521 499218 234587 499221
rect 234521 499216 235060 499218
rect 234521 499160 234526 499216
rect 234582 499160 235060 499216
rect 234521 499158 235060 499160
rect 234521 499155 234587 499158
rect 453941 498538 454007 498541
rect 451444 498536 454007 498538
rect 451444 498480 453946 498536
rect 454002 498480 454007 498536
rect 451444 498478 454007 498480
rect 453941 498475 454007 498478
rect 231526 497796 231532 497860
rect 231596 497858 231602 497860
rect 231596 497798 235060 497858
rect 583520 497844 584960 498084
rect 231596 497796 231602 497798
rect 454166 497178 454172 497180
rect 451444 497118 454172 497178
rect 454166 497116 454172 497118
rect 454236 497116 454242 497180
rect 232037 496498 232103 496501
rect 232037 496496 235060 496498
rect 232037 496440 232042 496496
rect 232098 496440 235060 496496
rect 232037 496438 235060 496440
rect 232037 496435 232103 496438
rect 233141 495138 233207 495141
rect 451733 495138 451799 495141
rect 233141 495136 235060 495138
rect 233141 495080 233146 495136
rect 233202 495080 235060 495136
rect 233141 495078 235060 495080
rect 451444 495136 451799 495138
rect 451444 495080 451738 495136
rect 451794 495080 451799 495136
rect 451444 495078 451799 495080
rect 233141 495075 233207 495078
rect 451733 495075 451799 495078
rect 232865 493778 232931 493781
rect 232865 493776 235060 493778
rect 232865 493720 232870 493776
rect 232926 493720 235060 493776
rect 232865 493718 235060 493720
rect 232865 493715 232931 493718
rect 451406 493716 451412 493780
rect 451476 493716 451482 493780
rect 453941 492418 454007 492421
rect 451444 492416 454007 492418
rect 228582 491268 228588 491332
rect 228652 491330 228658 491332
rect 235030 491330 235090 492388
rect 451444 492360 453946 492416
rect 454002 492360 454007 492416
rect 451444 492358 454007 492360
rect 453941 492355 454007 492358
rect 228652 491270 235090 491330
rect 228652 491268 228658 491270
rect 452653 491058 452719 491061
rect 451444 491056 452719 491058
rect 451444 491000 452658 491056
rect 452714 491000 452719 491056
rect 451444 490998 452719 491000
rect 452653 490995 452719 490998
rect 232037 489698 232103 489701
rect 453757 489698 453823 489701
rect 232037 489696 235060 489698
rect 232037 489640 232042 489696
rect 232098 489640 235060 489696
rect 232037 489638 235060 489640
rect 451444 489696 453823 489698
rect 451444 489640 453762 489696
rect 453818 489640 453823 489696
rect 451444 489638 453823 489640
rect 232037 489635 232103 489638
rect 453757 489635 453823 489638
rect -960 488596 480 488836
rect 453941 488338 454007 488341
rect 451444 488336 454007 488338
rect 451444 488280 453946 488336
rect 454002 488280 454007 488336
rect 451444 488278 454007 488280
rect 453941 488275 454007 488278
rect 231853 486978 231919 486981
rect 453757 486978 453823 486981
rect 231853 486976 235060 486978
rect 231853 486920 231858 486976
rect 231914 486920 235060 486976
rect 231853 486918 235060 486920
rect 451444 486976 453823 486978
rect 451444 486920 453762 486976
rect 453818 486920 453823 486976
rect 451444 486918 453823 486920
rect 231853 486915 231919 486918
rect 453757 486915 453823 486918
rect 232037 485618 232103 485621
rect 453941 485618 454007 485621
rect 232037 485616 235060 485618
rect 232037 485560 232042 485616
rect 232098 485560 235060 485616
rect 232037 485558 235060 485560
rect 451444 485616 454007 485618
rect 451444 485560 453946 485616
rect 454002 485560 454007 485616
rect 451444 485558 454007 485560
rect 232037 485555 232103 485558
rect 453941 485555 454007 485558
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 234153 484258 234219 484261
rect 459502 484258 459508 484260
rect 234153 484256 235060 484258
rect 234153 484200 234158 484256
rect 234214 484200 235060 484256
rect 234153 484198 235060 484200
rect 451444 484198 459508 484258
rect 234153 484195 234219 484198
rect 459502 484196 459508 484198
rect 459572 484196 459578 484260
rect 232037 482898 232103 482901
rect 453205 482898 453271 482901
rect 232037 482896 235060 482898
rect 232037 482840 232042 482896
rect 232098 482840 235060 482896
rect 232037 482838 235060 482840
rect 451444 482896 453271 482898
rect 451444 482840 453210 482896
rect 453266 482840 453271 482896
rect 451444 482838 453271 482840
rect 232037 482835 232103 482838
rect 453205 482835 453271 482838
rect 232037 481538 232103 481541
rect 453757 481538 453823 481541
rect 232037 481536 235060 481538
rect 232037 481480 232042 481536
rect 232098 481480 235060 481536
rect 232037 481478 235060 481480
rect 451444 481536 453823 481538
rect 451444 481480 453762 481536
rect 453818 481480 453823 481536
rect 451444 481478 453823 481480
rect 232037 481475 232103 481478
rect 453757 481475 453823 481478
rect 451825 480178 451891 480181
rect 451444 480176 451891 480178
rect 451444 480120 451830 480176
rect 451886 480120 451891 480176
rect 451444 480118 451891 480120
rect 451825 480115 451891 480118
rect 231393 479498 231459 479501
rect 231393 479496 235060 479498
rect 231393 479440 231398 479496
rect 231454 479440 235060 479496
rect 231393 479438 235060 479440
rect 231393 479435 231459 479438
rect 453757 478818 453823 478821
rect 451444 478816 453823 478818
rect 451444 478760 453762 478816
rect 453818 478760 453823 478816
rect 451444 478758 453823 478760
rect 453757 478755 453823 478758
rect 232037 478138 232103 478141
rect 232037 478136 235060 478138
rect 232037 478080 232042 478136
rect 232098 478080 235060 478136
rect 232037 478078 235060 478080
rect 232037 478075 232103 478078
rect 453849 477458 453915 477461
rect 451444 477456 453915 477458
rect 451444 477400 453854 477456
rect 453910 477400 453915 477456
rect 451444 477398 453915 477400
rect 453849 477395 453915 477398
rect 231301 476778 231367 476781
rect 231301 476776 235060 476778
rect 231301 476720 231306 476776
rect 231362 476720 235060 476776
rect 231301 476718 235060 476720
rect 231301 476715 231367 476718
rect 453941 476098 454007 476101
rect 451444 476096 454007 476098
rect 451444 476040 453946 476096
rect 454002 476040 454007 476096
rect 451444 476038 454007 476040
rect 453941 476035 454007 476038
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 232037 475418 232103 475421
rect 232037 475416 235060 475418
rect 232037 475360 232042 475416
rect 232098 475360 235060 475416
rect 232037 475358 235060 475360
rect 232037 475355 232103 475358
rect 231853 474058 231919 474061
rect 452101 474058 452167 474061
rect 231853 474056 235060 474058
rect 231853 474000 231858 474056
rect 231914 474000 235060 474056
rect 231853 473998 235060 474000
rect 451444 474056 452167 474058
rect 451444 474000 452106 474056
rect 452162 474000 452167 474056
rect 451444 473998 452167 474000
rect 231853 473995 231919 473998
rect 452101 473995 452167 473998
rect 232037 472698 232103 472701
rect 453941 472698 454007 472701
rect 232037 472696 235060 472698
rect 232037 472640 232042 472696
rect 232098 472640 235060 472696
rect 232037 472638 235060 472640
rect 451444 472696 454007 472698
rect 451444 472640 453946 472696
rect 454002 472640 454007 472696
rect 451444 472638 454007 472640
rect 232037 472635 232103 472638
rect 453941 472635 454007 472638
rect 579613 471474 579679 471477
rect 583520 471474 584960 471564
rect 579613 471472 584960 471474
rect 579613 471416 579618 471472
rect 579674 471416 584960 471472
rect 579613 471414 584960 471416
rect 579613 471411 579679 471414
rect 232037 471338 232103 471341
rect 453757 471338 453823 471341
rect 232037 471336 235060 471338
rect 232037 471280 232042 471336
rect 232098 471280 235060 471336
rect 232037 471278 235060 471280
rect 451444 471336 453823 471338
rect 451444 471280 453762 471336
rect 453818 471280 453823 471336
rect 583520 471324 584960 471414
rect 451444 471278 453823 471280
rect 232037 471275 232103 471278
rect 453757 471275 453823 471278
rect 233550 469916 233556 469980
rect 233620 469978 233626 469980
rect 453941 469978 454007 469981
rect 233620 469918 235060 469978
rect 451444 469976 454007 469978
rect 451444 469920 453946 469976
rect 454002 469920 454007 469976
rect 451444 469918 454007 469920
rect 233620 469916 233626 469918
rect 453941 469915 454007 469918
rect 234245 468618 234311 468621
rect 452653 468618 452719 468621
rect 234245 468616 235060 468618
rect 234245 468560 234250 468616
rect 234306 468560 235060 468616
rect 234245 468558 235060 468560
rect 451444 468616 452719 468618
rect 451444 468560 452658 468616
rect 452714 468560 452719 468616
rect 451444 468558 452719 468560
rect 234245 468555 234311 468558
rect 452653 468555 452719 468558
rect 232998 467196 233004 467260
rect 233068 467258 233074 467260
rect 453573 467258 453639 467261
rect 233068 467198 235060 467258
rect 451444 467256 453639 467258
rect 451444 467200 453578 467256
rect 453634 467200 453639 467256
rect 451444 467198 453639 467200
rect 233068 467196 233074 467198
rect 453573 467195 453639 467198
rect 232037 465898 232103 465901
rect 454217 465898 454283 465901
rect 232037 465896 235060 465898
rect 232037 465840 232042 465896
rect 232098 465840 235060 465896
rect 232037 465838 235060 465840
rect 451444 465896 454283 465898
rect 451444 465840 454222 465896
rect 454278 465840 454283 465896
rect 451444 465838 454283 465840
rect 232037 465835 232103 465838
rect 454217 465835 454283 465838
rect 232037 464538 232103 464541
rect 453205 464538 453271 464541
rect 232037 464536 235060 464538
rect 232037 464480 232042 464536
rect 232098 464480 235060 464536
rect 232037 464478 235060 464480
rect 451444 464536 453271 464538
rect 451444 464480 453210 464536
rect 453266 464480 453271 464536
rect 451444 464478 453271 464480
rect 232037 464475 232103 464478
rect 453205 464475 453271 464478
rect 232037 463178 232103 463181
rect 453941 463178 454007 463181
rect 232037 463176 235060 463178
rect 232037 463120 232042 463176
rect 232098 463120 235060 463176
rect 232037 463118 235060 463120
rect 451444 463176 454007 463178
rect 451444 463120 453946 463176
rect 454002 463120 454007 463176
rect 451444 463118 454007 463120
rect 232037 463115 232103 463118
rect 453941 463115 454007 463118
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 232037 461818 232103 461821
rect 455454 461818 455460 461820
rect 232037 461816 235060 461818
rect 232037 461760 232042 461816
rect 232098 461760 235060 461816
rect 232037 461758 235060 461760
rect 451444 461758 455460 461818
rect 232037 461755 232103 461758
rect 455454 461756 455460 461758
rect 455524 461756 455530 461820
rect 232037 460458 232103 460461
rect 453941 460458 454007 460461
rect 232037 460456 235060 460458
rect 232037 460400 232042 460456
rect 232098 460400 235060 460456
rect 232037 460398 235060 460400
rect 451444 460456 454007 460458
rect 451444 460400 453946 460456
rect 454002 460400 454007 460456
rect 451444 460398 454007 460400
rect 232037 460395 232103 460398
rect 453941 460395 454007 460398
rect 452653 459098 452719 459101
rect 451444 459096 452719 459098
rect 451444 459040 452658 459096
rect 452714 459040 452719 459096
rect 451444 459038 452719 459040
rect 452653 459035 452719 459038
rect 231945 458418 232011 458421
rect 231945 458416 235060 458418
rect 231945 458360 231950 458416
rect 232006 458360 235060 458416
rect 231945 458358 235060 458360
rect 231945 458355 232011 458358
rect 580533 458146 580599 458149
rect 583520 458146 584960 458236
rect 580533 458144 584960 458146
rect 580533 458088 580538 458144
rect 580594 458088 584960 458144
rect 580533 458086 584960 458088
rect 580533 458083 580599 458086
rect 583520 457996 584960 458086
rect 452009 457738 452075 457741
rect 451444 457736 452075 457738
rect 451444 457680 452014 457736
rect 452070 457680 452075 457736
rect 451444 457678 452075 457680
rect 452009 457675 452075 457678
rect 232037 457058 232103 457061
rect 232037 457056 235060 457058
rect 232037 457000 232042 457056
rect 232098 457000 235060 457056
rect 232037 456998 235060 457000
rect 232037 456995 232103 456998
rect 453665 456378 453731 456381
rect 451444 456376 453731 456378
rect 451444 456320 453670 456376
rect 453726 456320 453731 456376
rect 451444 456318 453731 456320
rect 453665 456315 453731 456318
rect 231945 455698 232011 455701
rect 231945 455696 235060 455698
rect 231945 455640 231950 455696
rect 232006 455640 235060 455696
rect 231945 455638 235060 455640
rect 231945 455635 232011 455638
rect 232037 454338 232103 454341
rect 453941 454338 454007 454341
rect 232037 454336 235060 454338
rect 232037 454280 232042 454336
rect 232098 454280 235060 454336
rect 232037 454278 235060 454280
rect 451444 454336 454007 454338
rect 451444 454280 453946 454336
rect 454002 454280 454007 454336
rect 451444 454278 454007 454280
rect 232037 454275 232103 454278
rect 453941 454275 454007 454278
rect 232037 452978 232103 452981
rect 453941 452978 454007 452981
rect 232037 452976 235060 452978
rect 232037 452920 232042 452976
rect 232098 452920 235060 452976
rect 232037 452918 235060 452920
rect 451444 452976 454007 452978
rect 451444 452920 453946 452976
rect 454002 452920 454007 452976
rect 451444 452918 454007 452920
rect 232037 452915 232103 452918
rect 453941 452915 454007 452918
rect 232037 451618 232103 451621
rect 453021 451618 453087 451621
rect 232037 451616 235060 451618
rect 232037 451560 232042 451616
rect 232098 451560 235060 451616
rect 232037 451558 235060 451560
rect 451444 451616 453087 451618
rect 451444 451560 453026 451616
rect 453082 451560 453087 451616
rect 451444 451558 453087 451560
rect 232037 451555 232103 451558
rect 453021 451555 453087 451558
rect 232865 450258 232931 450261
rect 453573 450258 453639 450261
rect 232865 450256 235060 450258
rect 232865 450200 232870 450256
rect 232926 450200 235060 450256
rect 232865 450198 235060 450200
rect 451444 450256 453639 450258
rect 451444 450200 453578 450256
rect 453634 450200 453639 450256
rect 451444 450198 453639 450200
rect 232865 450195 232931 450198
rect 453573 450195 453639 450198
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 231485 448898 231551 448901
rect 454350 448898 454356 448900
rect 231485 448896 235060 448898
rect 231485 448840 231490 448896
rect 231546 448840 235060 448896
rect 231485 448838 235060 448840
rect 451444 448838 454356 448898
rect 231485 448835 231551 448838
rect 454350 448836 454356 448838
rect 454420 448836 454426 448900
rect 233182 447476 233188 447540
rect 233252 447538 233258 447540
rect 453021 447538 453087 447541
rect 233252 447478 235060 447538
rect 451444 447536 453087 447538
rect 451444 447480 453026 447536
rect 453082 447480 453087 447536
rect 451444 447478 453087 447480
rect 233252 447476 233258 447478
rect 453021 447475 453087 447478
rect 454166 446178 454172 446180
rect 451444 446118 454172 446178
rect 454166 446116 454172 446118
rect 454236 446116 454242 446180
rect 232313 444818 232379 444821
rect 453941 444818 454007 444821
rect 232313 444816 235060 444818
rect 232313 444760 232318 444816
rect 232374 444760 235060 444816
rect 232313 444758 235060 444760
rect 451444 444816 454007 444818
rect 451444 444760 453946 444816
rect 454002 444760 454007 444816
rect 451444 444758 454007 444760
rect 232313 444755 232379 444758
rect 453941 444755 454007 444758
rect 583520 444668 584960 444908
rect 232037 443458 232103 443461
rect 457110 443458 457116 443460
rect 232037 443456 235060 443458
rect 232037 443400 232042 443456
rect 232098 443400 235060 443456
rect 232037 443398 235060 443400
rect 451444 443398 457116 443458
rect 232037 443395 232103 443398
rect 457110 443396 457116 443398
rect 457180 443396 457186 443460
rect 232037 442098 232103 442101
rect 232037 442096 235060 442098
rect 232037 442040 232042 442096
rect 232098 442040 235060 442096
rect 232037 442038 235060 442040
rect 232037 442035 232103 442038
rect 451414 441690 451474 442068
rect 462262 441690 462268 441692
rect 451414 441630 462268 441690
rect 462262 441628 462268 441630
rect 462332 441628 462338 441692
rect 232037 440738 232103 440741
rect 453941 440738 454007 440741
rect 232037 440736 235060 440738
rect 232037 440680 232042 440736
rect 232098 440680 235060 440736
rect 232037 440678 235060 440680
rect 451444 440736 454007 440738
rect 451444 440680 453946 440736
rect 454002 440680 454007 440736
rect 451444 440678 454007 440680
rect 232037 440675 232103 440678
rect 453941 440675 454007 440678
rect 453849 439378 453915 439381
rect 451444 439376 453915 439378
rect 451444 439320 453854 439376
rect 453910 439320 453915 439376
rect 451444 439318 453915 439320
rect 453849 439315 453915 439318
rect 234245 438698 234311 438701
rect 234245 438696 235060 438698
rect 234245 438640 234250 438696
rect 234306 438640 235060 438696
rect 234245 438638 235060 438640
rect 234245 438635 234311 438638
rect 453941 438018 454007 438021
rect 451444 438016 454007 438018
rect 451444 437960 453946 438016
rect 454002 437960 454007 438016
rect 451444 437958 454007 437960
rect 453941 437955 454007 437958
rect 232814 437276 232820 437340
rect 232884 437338 232890 437340
rect 232884 437278 235060 437338
rect 232884 437276 232890 437278
rect -960 436508 480 436748
rect 453941 436658 454007 436661
rect 451444 436656 454007 436658
rect 451444 436600 453946 436656
rect 454002 436600 454007 436656
rect 451444 436598 454007 436600
rect 453941 436595 454007 436598
rect 232589 435978 232655 435981
rect 232589 435976 235060 435978
rect 232589 435920 232594 435976
rect 232650 435920 235060 435976
rect 232589 435918 235060 435920
rect 232589 435915 232655 435918
rect 453665 435298 453731 435301
rect 451444 435296 453731 435298
rect 451444 435240 453670 435296
rect 453726 435240 453731 435296
rect 451444 435238 453731 435240
rect 453665 435235 453731 435238
rect 231945 434618 232011 434621
rect 231945 434616 235060 434618
rect 231945 434560 231950 434616
rect 232006 434560 235060 434616
rect 231945 434558 235060 434560
rect 231945 434555 232011 434558
rect 232037 433258 232103 433261
rect 457294 433258 457300 433260
rect 232037 433256 235060 433258
rect 232037 433200 232042 433256
rect 232098 433200 235060 433256
rect 232037 433198 235060 433200
rect 451444 433198 457300 433258
rect 232037 433195 232103 433198
rect 457294 433196 457300 433198
rect 457364 433196 457370 433260
rect 231209 431898 231275 431901
rect 453941 431898 454007 431901
rect 231209 431896 235060 431898
rect 231209 431840 231214 431896
rect 231270 431840 235060 431896
rect 231209 431838 235060 431840
rect 451444 431896 454007 431898
rect 451444 431840 453946 431896
rect 454002 431840 454007 431896
rect 451444 431838 454007 431840
rect 231209 431835 231275 431838
rect 453941 431835 454007 431838
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 231853 430538 231919 430541
rect 452745 430538 452811 430541
rect 231853 430536 235060 430538
rect 231853 430480 231858 430536
rect 231914 430480 235060 430536
rect 231853 430478 235060 430480
rect 451444 430536 452811 430538
rect 451444 430480 452750 430536
rect 452806 430480 452811 430536
rect 451444 430478 452811 430480
rect 231853 430475 231919 430478
rect 452745 430475 452811 430478
rect 232037 429178 232103 429181
rect 453941 429178 454007 429181
rect 232037 429176 235060 429178
rect 232037 429120 232042 429176
rect 232098 429120 235060 429176
rect 232037 429118 235060 429120
rect 451444 429176 454007 429178
rect 451444 429120 453946 429176
rect 454002 429120 454007 429176
rect 451444 429118 454007 429120
rect 232037 429115 232103 429118
rect 453941 429115 454007 429118
rect 235022 427756 235028 427820
rect 235092 427756 235098 427820
rect 453021 427818 453087 427821
rect 451444 427816 453087 427818
rect 451444 427760 453026 427816
rect 453082 427760 453087 427816
rect 451444 427758 453087 427760
rect 453021 427755 453087 427758
rect 232037 426458 232103 426461
rect 453941 426458 454007 426461
rect 232037 426456 235060 426458
rect 232037 426400 232042 426456
rect 232098 426400 235060 426456
rect 232037 426398 235060 426400
rect 451444 426456 454007 426458
rect 451444 426400 453946 426456
rect 454002 426400 454007 426456
rect 451444 426398 454007 426400
rect 232037 426395 232103 426398
rect 453941 426395 454007 426398
rect 232037 425098 232103 425101
rect 453941 425098 454007 425101
rect 232037 425096 235060 425098
rect 232037 425040 232042 425096
rect 232098 425040 235060 425096
rect 232037 425038 235060 425040
rect 451444 425096 454007 425098
rect 451444 425040 453946 425096
rect 454002 425040 454007 425096
rect 451444 425038 454007 425040
rect 232037 425035 232103 425038
rect 453941 425035 454007 425038
rect 232037 423738 232103 423741
rect 452745 423738 452811 423741
rect 232037 423736 235060 423738
rect -960 423602 480 423692
rect 232037 423680 232042 423736
rect 232098 423680 235060 423736
rect 232037 423678 235060 423680
rect 451444 423736 452811 423738
rect 451444 423680 452750 423736
rect 452806 423680 452811 423736
rect 451444 423678 452811 423680
rect 232037 423675 232103 423678
rect 452745 423675 452811 423678
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 232773 422378 232839 422381
rect 454534 422378 454540 422380
rect 232773 422376 235060 422378
rect 232773 422320 232778 422376
rect 232834 422320 235060 422376
rect 232773 422318 235060 422320
rect 451444 422318 454540 422378
rect 232773 422315 232839 422318
rect 454534 422316 454540 422318
rect 454604 422316 454610 422380
rect 234061 421018 234127 421021
rect 453941 421018 454007 421021
rect 234061 421016 235060 421018
rect 234061 420960 234066 421016
rect 234122 420960 235060 421016
rect 234061 420958 235060 420960
rect 451444 421016 454007 421018
rect 451444 420960 453946 421016
rect 454002 420960 454007 421016
rect 451444 420958 454007 420960
rect 234061 420955 234127 420958
rect 453941 420955 454007 420958
rect 232037 419658 232103 419661
rect 232037 419656 235060 419658
rect 232037 419600 232042 419656
rect 232098 419600 235060 419656
rect 232037 419598 235060 419600
rect 232037 419595 232103 419598
rect 453665 418298 453731 418301
rect 451444 418296 453731 418298
rect 451444 418240 453670 418296
rect 453726 418240 453731 418296
rect 451444 418238 453731 418240
rect 453665 418235 453731 418238
rect 579705 418298 579771 418301
rect 583520 418298 584960 418388
rect 579705 418296 584960 418298
rect 579705 418240 579710 418296
rect 579766 418240 584960 418296
rect 579705 418238 584960 418240
rect 579705 418235 579771 418238
rect 583520 418148 584960 418238
rect 234705 417618 234771 417621
rect 234705 417616 235060 417618
rect 234705 417560 234710 417616
rect 234766 417560 235060 417616
rect 234705 417558 235060 417560
rect 234705 417555 234771 417558
rect 453205 416938 453271 416941
rect 451444 416936 453271 416938
rect 451444 416880 453210 416936
rect 453266 416880 453271 416936
rect 451444 416878 453271 416880
rect 453205 416875 453271 416878
rect 231945 416258 232011 416261
rect 231945 416256 235060 416258
rect 231945 416200 231950 416256
rect 232006 416200 235060 416256
rect 231945 416198 235060 416200
rect 231945 416195 232011 416198
rect 456006 415578 456012 415580
rect 451444 415518 456012 415578
rect 456006 415516 456012 415518
rect 456076 415516 456082 415580
rect 229870 414836 229876 414900
rect 229940 414898 229946 414900
rect 229940 414838 235060 414898
rect 229940 414836 229946 414838
rect 232037 413538 232103 413541
rect 453941 413538 454007 413541
rect 232037 413536 235060 413538
rect 232037 413480 232042 413536
rect 232098 413480 235060 413536
rect 232037 413478 235060 413480
rect 451444 413536 454007 413538
rect 451444 413480 453946 413536
rect 454002 413480 454007 413536
rect 451444 413478 454007 413480
rect 232037 413475 232103 413478
rect 453941 413475 454007 413478
rect 233049 412178 233115 412181
rect 455822 412178 455828 412180
rect 233049 412176 235060 412178
rect 233049 412120 233054 412176
rect 233110 412120 235060 412176
rect 233049 412118 235060 412120
rect 451444 412118 455828 412178
rect 233049 412115 233115 412118
rect 455822 412116 455828 412118
rect 455892 412116 455898 412180
rect 232037 410818 232103 410821
rect 452694 410818 452700 410820
rect 232037 410816 235060 410818
rect 232037 410760 232042 410816
rect 232098 410760 235060 410816
rect 232037 410758 235060 410760
rect 451444 410758 452700 410818
rect 232037 410755 232103 410758
rect 452694 410756 452700 410758
rect 452764 410756 452770 410820
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 451958 409940 451964 410004
rect 452028 410002 452034 410004
rect 452837 410002 452903 410005
rect 452028 410000 452903 410002
rect 452028 409944 452842 410000
rect 452898 409944 452903 410000
rect 452028 409942 452903 409944
rect 452028 409940 452034 409942
rect 452837 409939 452903 409942
rect 234337 409458 234403 409461
rect 452653 409458 452719 409461
rect 234337 409456 235060 409458
rect 234337 409400 234342 409456
rect 234398 409400 235060 409456
rect 234337 409398 235060 409400
rect 451444 409456 452719 409458
rect 451444 409400 452658 409456
rect 452714 409400 452719 409456
rect 451444 409398 452719 409400
rect 234337 409395 234403 409398
rect 452653 409395 452719 409398
rect 232037 408098 232103 408101
rect 453757 408098 453823 408101
rect 232037 408096 235060 408098
rect 232037 408040 232042 408096
rect 232098 408040 235060 408096
rect 232037 408038 235060 408040
rect 451444 408096 453823 408098
rect 451444 408040 453762 408096
rect 453818 408040 453823 408096
rect 451444 408038 453823 408040
rect 232037 408035 232103 408038
rect 453757 408035 453823 408038
rect 232630 406676 232636 406740
rect 232700 406738 232706 406740
rect 453941 406738 454007 406741
rect 232700 406678 235060 406738
rect 451444 406736 454007 406738
rect 451444 406680 453946 406736
rect 454002 406680 454007 406736
rect 451444 406678 454007 406680
rect 232700 406676 232706 406678
rect 453941 406675 454007 406678
rect 234337 405378 234403 405381
rect 453757 405378 453823 405381
rect 234337 405376 235060 405378
rect 234337 405320 234342 405376
rect 234398 405320 235060 405376
rect 234337 405318 235060 405320
rect 451444 405376 453823 405378
rect 451444 405320 453762 405376
rect 453818 405320 453823 405376
rect 451444 405318 453823 405320
rect 234337 405315 234403 405318
rect 453757 405315 453823 405318
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 232405 404018 232471 404021
rect 232405 404016 235060 404018
rect 232405 403960 232410 404016
rect 232466 403960 235060 404016
rect 232405 403958 235060 403960
rect 232405 403955 232471 403958
rect 450854 403956 450860 404020
rect 450924 403956 450930 404020
rect 232037 402658 232103 402661
rect 453941 402658 454007 402661
rect 232037 402656 235060 402658
rect 232037 402600 232042 402656
rect 232098 402600 235060 402656
rect 232037 402598 235060 402600
rect 451444 402656 454007 402658
rect 451444 402600 453946 402656
rect 454002 402600 454007 402656
rect 451444 402598 454007 402600
rect 232037 402595 232103 402598
rect 453941 402595 454007 402598
rect 234153 401298 234219 401301
rect 452653 401298 452719 401301
rect 234153 401296 235060 401298
rect 234153 401240 234158 401296
rect 234214 401240 235060 401296
rect 234153 401238 235060 401240
rect 451444 401296 452719 401298
rect 451444 401240 452658 401296
rect 452714 401240 452719 401296
rect 451444 401238 452719 401240
rect 234153 401235 234219 401238
rect 452653 401235 452719 401238
rect 232037 399938 232103 399941
rect 453757 399938 453823 399941
rect 232037 399936 235060 399938
rect 232037 399880 232042 399936
rect 232098 399880 235060 399936
rect 232037 399878 235060 399880
rect 451444 399936 453823 399938
rect 451444 399880 453762 399936
rect 453818 399880 453823 399936
rect 451444 399878 453823 399880
rect 232037 399875 232103 399878
rect 453757 399875 453823 399878
rect 453062 398578 453068 398580
rect 451444 398518 453068 398578
rect 453062 398516 453068 398518
rect 453132 398516 453138 398580
rect 232037 397898 232103 397901
rect 232037 397896 235060 397898
rect 232037 397840 232042 397896
rect 232098 397840 235060 397896
rect 232037 397838 235060 397840
rect 232037 397835 232103 397838
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 231945 396538 232011 396541
rect 231945 396536 235060 396538
rect 231945 396480 231950 396536
rect 232006 396480 235060 396536
rect 231945 396478 235060 396480
rect 231945 396475 232011 396478
rect 453757 395858 453823 395861
rect 451444 395856 453823 395858
rect 451444 395800 453762 395856
rect 453818 395800 453823 395856
rect 451444 395798 453823 395800
rect 453757 395795 453823 395798
rect 232037 395178 232103 395181
rect 232037 395176 235060 395178
rect 232037 395120 232042 395176
rect 232098 395120 235060 395176
rect 232037 395118 235060 395120
rect 232037 395115 232103 395118
rect 453757 394498 453823 394501
rect 451444 394496 453823 394498
rect 451444 394440 453762 394496
rect 453818 394440 453823 394496
rect 451444 394438 453823 394440
rect 453757 394435 453823 394438
rect 232405 393818 232471 393821
rect 232405 393816 235060 393818
rect 232405 393760 232410 393816
rect 232466 393760 235060 393816
rect 232405 393758 235060 393760
rect 232405 393755 232471 393758
rect 233969 392458 234035 392461
rect 453941 392458 454007 392461
rect 233969 392456 235060 392458
rect 233969 392400 233974 392456
rect 234030 392400 235060 392456
rect 233969 392398 235060 392400
rect 451444 392456 454007 392458
rect 451444 392400 453946 392456
rect 454002 392400 454007 392456
rect 451444 392398 454007 392400
rect 233969 392395 234035 392398
rect 453941 392395 454007 392398
rect 583520 391628 584960 391868
rect 232037 391098 232103 391101
rect 452193 391098 452259 391101
rect 232037 391096 235060 391098
rect 232037 391040 232042 391096
rect 232098 391040 235060 391096
rect 232037 391038 235060 391040
rect 451444 391096 452259 391098
rect 451444 391040 452198 391096
rect 452254 391040 452259 391096
rect 451444 391038 452259 391040
rect 232037 391035 232103 391038
rect 452193 391035 452259 391038
rect 231117 389738 231183 389741
rect 453941 389738 454007 389741
rect 231117 389736 235060 389738
rect 231117 389680 231122 389736
rect 231178 389680 235060 389736
rect 231117 389678 235060 389680
rect 451444 389736 454007 389738
rect 451444 389680 453946 389736
rect 454002 389680 454007 389736
rect 451444 389678 454007 389680
rect 231117 389675 231183 389678
rect 453941 389675 454007 389678
rect 232446 388316 232452 388380
rect 232516 388378 232522 388380
rect 452837 388378 452903 388381
rect 232516 388318 235060 388378
rect 451444 388376 452903 388378
rect 451444 388320 452842 388376
rect 452898 388320 452903 388376
rect 451444 388318 452903 388320
rect 232516 388316 232522 388318
rect 452837 388315 452903 388318
rect 235206 386956 235212 387020
rect 235276 386956 235282 387020
rect 453941 387018 454007 387021
rect 451444 387016 454007 387018
rect 451444 386960 453946 387016
rect 454002 386960 454007 387016
rect 451444 386958 454007 386960
rect 453941 386955 454007 386958
rect 232037 385658 232103 385661
rect 453941 385658 454007 385661
rect 232037 385656 235060 385658
rect 232037 385600 232042 385656
rect 232098 385600 235060 385656
rect 232037 385598 235060 385600
rect 451444 385656 454007 385658
rect 451444 385600 453946 385656
rect 454002 385600 454007 385656
rect 451444 385598 454007 385600
rect 232037 385595 232103 385598
rect 453941 385595 454007 385598
rect -960 384284 480 384524
rect 232037 384298 232103 384301
rect 453941 384298 454007 384301
rect 232037 384296 235060 384298
rect 232037 384240 232042 384296
rect 232098 384240 235060 384296
rect 232037 384238 235060 384240
rect 451444 384296 454007 384298
rect 451444 384240 453946 384296
rect 454002 384240 454007 384296
rect 451444 384238 454007 384240
rect 232037 384235 232103 384238
rect 453941 384235 454007 384238
rect 232681 382938 232747 382941
rect 453205 382938 453271 382941
rect 232681 382936 235060 382938
rect 232681 382880 232686 382936
rect 232742 382880 235060 382936
rect 232681 382878 235060 382880
rect 451444 382936 453271 382938
rect 451444 382880 453210 382936
rect 453266 382880 453271 382936
rect 451444 382878 453271 382880
rect 232681 382875 232747 382878
rect 453205 382875 453271 382878
rect 233785 380218 233851 380221
rect 453113 380218 453179 380221
rect 233785 380216 235060 380218
rect 233785 380160 233790 380216
rect 233846 380160 235060 380216
rect 233785 380158 235060 380160
rect 451444 380216 453179 380218
rect 451444 380160 453118 380216
rect 453174 380160 453179 380216
rect 451444 380158 453179 380160
rect 233785 380155 233851 380158
rect 453113 380155 453179 380158
rect 232037 378858 232103 378861
rect 453757 378858 453823 378861
rect 232037 378856 235060 378858
rect 232037 378800 232042 378856
rect 232098 378800 235060 378856
rect 232037 378798 235060 378800
rect 451444 378856 453823 378858
rect 451444 378800 453762 378856
rect 453818 378800 453823 378856
rect 451444 378798 453823 378800
rect 232037 378795 232103 378798
rect 453757 378795 453823 378798
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 232129 376818 232195 376821
rect 232129 376816 235060 376818
rect 232129 376760 232134 376816
rect 232190 376760 235060 376816
rect 232129 376758 235060 376760
rect 232129 376755 232195 376758
rect 453757 376138 453823 376141
rect 451444 376136 453823 376138
rect 451444 376080 453762 376136
rect 453818 376080 453823 376136
rect 451444 376078 453823 376080
rect 453757 376075 453823 376078
rect 232037 375458 232103 375461
rect 232037 375456 235060 375458
rect 232037 375400 232042 375456
rect 232098 375400 235060 375456
rect 232037 375398 235060 375400
rect 232037 375395 232103 375398
rect 452745 374778 452811 374781
rect 451444 374776 452811 374778
rect 451444 374720 452750 374776
rect 452806 374720 452811 374776
rect 451444 374718 452811 374720
rect 452745 374715 452811 374718
rect 231853 374098 231919 374101
rect 231853 374096 235060 374098
rect 231853 374040 231858 374096
rect 231914 374040 235060 374096
rect 231853 374038 235060 374040
rect 231853 374035 231919 374038
rect 232037 372738 232103 372741
rect 453941 372738 454007 372741
rect 232037 372736 235060 372738
rect 232037 372680 232042 372736
rect 232098 372680 235060 372736
rect 232037 372678 235060 372680
rect 451444 372736 454007 372738
rect 451444 372680 453946 372736
rect 454002 372680 454007 372736
rect 451444 372678 454007 372680
rect 232037 372675 232103 372678
rect 453941 372675 454007 372678
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 232037 371378 232103 371381
rect 453757 371378 453823 371381
rect 232037 371376 235060 371378
rect 232037 371320 232042 371376
rect 232098 371320 235060 371376
rect 232037 371318 235060 371320
rect 451444 371376 453823 371378
rect 451444 371320 453762 371376
rect 453818 371320 453823 371376
rect 451444 371318 453823 371320
rect 232037 371315 232103 371318
rect 453757 371315 453823 371318
rect 234797 370018 234863 370021
rect 453757 370018 453823 370021
rect 234797 370016 235060 370018
rect 234797 369960 234802 370016
rect 234858 369960 235060 370016
rect 234797 369958 235060 369960
rect 451444 370016 453823 370018
rect 451444 369960 453762 370016
rect 453818 369960 453823 370016
rect 451444 369958 453823 369960
rect 234797 369955 234863 369958
rect 453757 369955 453823 369958
rect 232037 368658 232103 368661
rect 453757 368658 453823 368661
rect 232037 368656 235060 368658
rect 232037 368600 232042 368656
rect 232098 368600 235060 368656
rect 232037 368598 235060 368600
rect 451444 368656 453823 368658
rect 451444 368600 453762 368656
rect 453818 368600 453823 368656
rect 451444 368598 453823 368600
rect 232037 368595 232103 368598
rect 453757 368595 453823 368598
rect 231853 367298 231919 367301
rect 453941 367298 454007 367301
rect 231853 367296 235060 367298
rect 231853 367240 231858 367296
rect 231914 367240 235060 367296
rect 231853 367238 235060 367240
rect 451444 367296 454007 367298
rect 451444 367240 453946 367296
rect 454002 367240 454007 367296
rect 451444 367238 454007 367240
rect 231853 367235 231919 367238
rect 453941 367235 454007 367238
rect 453941 365938 454007 365941
rect 451444 365936 454007 365938
rect 451444 365880 453946 365936
rect 454002 365880 454007 365936
rect 451444 365878 454007 365880
rect 453941 365875 454007 365878
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 232497 364578 232563 364581
rect 453757 364578 453823 364581
rect 232497 364576 235060 364578
rect 232497 364520 232502 364576
rect 232558 364520 235060 364576
rect 232497 364518 235060 364520
rect 451444 364576 453823 364578
rect 451444 364520 453762 364576
rect 453818 364520 453823 364576
rect 451444 364518 453823 364520
rect 232497 364515 232563 364518
rect 453757 364515 453823 364518
rect 232037 363218 232103 363221
rect 453757 363218 453823 363221
rect 232037 363216 235060 363218
rect 232037 363160 232042 363216
rect 232098 363160 235060 363216
rect 232037 363158 235060 363160
rect 451444 363216 453823 363218
rect 451444 363160 453762 363216
rect 453818 363160 453823 363216
rect 451444 363158 453823 363160
rect 232037 363155 232103 363158
rect 453757 363155 453823 363158
rect 232037 361858 232103 361861
rect 453941 361858 454007 361861
rect 232037 361856 235060 361858
rect 232037 361800 232042 361856
rect 232098 361800 235060 361856
rect 232037 361798 235060 361800
rect 451444 361856 454007 361858
rect 451444 361800 453946 361856
rect 454002 361800 454007 361856
rect 451444 361798 454007 361800
rect 232037 361795 232103 361798
rect 453941 361795 454007 361798
rect 233877 360498 233943 360501
rect 233877 360496 235060 360498
rect 233877 360440 233882 360496
rect 233938 360440 235060 360496
rect 233877 360438 235060 360440
rect 233877 360435 233943 360438
rect 451414 360226 451474 360468
rect 460974 360226 460980 360228
rect 451414 360166 460980 360226
rect 460974 360164 460980 360166
rect 461044 360164 461050 360228
rect 233601 359138 233667 359141
rect 453941 359138 454007 359141
rect 233601 359136 235060 359138
rect 233601 359080 233606 359136
rect 233662 359080 235060 359136
rect 233601 359078 235060 359080
rect 451444 359136 454007 359138
rect 451444 359080 453946 359136
rect 454002 359080 454007 359136
rect 451444 359078 454007 359080
rect 233601 359075 233667 359078
rect 453941 359075 454007 359078
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 234429 358458 234495 358461
rect 235390 358458 235396 358460
rect 234429 358456 235396 358458
rect 234429 358400 234434 358456
rect 234490 358400 235396 358456
rect 234429 358398 235396 358400
rect 234429 358395 234495 358398
rect 235390 358396 235396 358398
rect 235460 358396 235466 358460
rect 453941 357778 454007 357781
rect 451444 357776 454007 357778
rect 451444 357720 453946 357776
rect 454002 357720 454007 357776
rect 451444 357718 454007 357720
rect 453941 357715 454007 357718
rect 232037 357098 232103 357101
rect 232037 357096 235060 357098
rect 232037 357040 232042 357096
rect 232098 357040 235060 357096
rect 232037 357038 235060 357040
rect 232037 357035 232103 357038
rect 453573 356418 453639 356421
rect 451444 356416 453639 356418
rect 451444 356360 453578 356416
rect 453634 356360 453639 356416
rect 451444 356358 453639 356360
rect 453573 356355 453639 356358
rect 233693 355738 233759 355741
rect 233693 355736 235060 355738
rect 233693 355680 233698 355736
rect 233754 355680 235060 355736
rect 233693 355678 235060 355680
rect 233693 355675 233759 355678
rect 452653 355058 452719 355061
rect 451444 355056 452719 355058
rect 451444 355000 452658 355056
rect 452714 355000 452719 355056
rect 451444 354998 452719 355000
rect 452653 354995 452719 354998
rect 232313 354378 232379 354381
rect 232313 354376 235060 354378
rect 232313 354320 232318 354376
rect 232374 354320 235060 354376
rect 232313 354318 235060 354320
rect 232313 354315 232379 354318
rect 453481 353698 453547 353701
rect 451444 353696 453547 353698
rect 451444 353640 453486 353696
rect 453542 353640 453547 353696
rect 451444 353638 453547 353640
rect 453481 353635 453547 353638
rect 232037 353018 232103 353021
rect 232037 353016 235060 353018
rect 232037 352960 232042 353016
rect 232098 352960 235060 353016
rect 232037 352958 235060 352960
rect 232037 352955 232103 352958
rect 580625 351930 580691 351933
rect 583520 351930 584960 352020
rect 580625 351928 584960 351930
rect 580625 351872 580630 351928
rect 580686 351872 584960 351928
rect 580625 351870 584960 351872
rect 580625 351867 580691 351870
rect 583520 351780 584960 351870
rect 232037 351658 232103 351661
rect 453246 351658 453252 351660
rect 232037 351656 235060 351658
rect 232037 351600 232042 351656
rect 232098 351600 235060 351656
rect 232037 351598 235060 351600
rect 451444 351598 453252 351658
rect 232037 351595 232103 351598
rect 453246 351596 453252 351598
rect 453316 351596 453322 351660
rect 232037 350298 232103 350301
rect 453665 350298 453731 350301
rect 232037 350296 235060 350298
rect 232037 350240 232042 350296
rect 232098 350240 235060 350296
rect 232037 350238 235060 350240
rect 451444 350296 453731 350298
rect 451444 350240 453670 350296
rect 453726 350240 453731 350296
rect 451444 350238 453731 350240
rect 232037 350235 232103 350238
rect 453665 350235 453731 350238
rect 232037 348938 232103 348941
rect 453941 348938 454007 348941
rect 232037 348936 235060 348938
rect 232037 348880 232042 348936
rect 232098 348880 235060 348936
rect 232037 348878 235060 348880
rect 451444 348936 454007 348938
rect 451444 348880 453946 348936
rect 454002 348880 454007 348936
rect 451444 348878 454007 348880
rect 232037 348875 232103 348878
rect 453941 348875 454007 348878
rect 232589 347578 232655 347581
rect 453941 347578 454007 347581
rect 232589 347576 235060 347578
rect 232589 347520 232594 347576
rect 232650 347520 235060 347576
rect 232589 347518 235060 347520
rect 451444 347576 454007 347578
rect 451444 347520 453946 347576
rect 454002 347520 454007 347576
rect 451444 347518 454007 347520
rect 232589 347515 232655 347518
rect 453941 347515 454007 347518
rect 232037 346218 232103 346221
rect 453205 346218 453271 346221
rect 232037 346216 235060 346218
rect 232037 346160 232042 346216
rect 232098 346160 235060 346216
rect 232037 346158 235060 346160
rect 451444 346216 453271 346218
rect 451444 346160 453210 346216
rect 453266 346160 453271 346216
rect 451444 346158 453271 346160
rect 232037 346155 232103 346158
rect 453205 346155 453271 346158
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 231945 344858 232011 344861
rect 452929 344858 452995 344861
rect 231945 344856 235060 344858
rect 231945 344800 231950 344856
rect 232006 344800 235060 344856
rect 231945 344798 235060 344800
rect 451444 344856 452995 344858
rect 451444 344800 452934 344856
rect 452990 344800 452995 344856
rect 451444 344798 452995 344800
rect 231945 344795 232011 344798
rect 452929 344795 452995 344798
rect 232037 343498 232103 343501
rect 453941 343498 454007 343501
rect 232037 343496 235060 343498
rect 232037 343440 232042 343496
rect 232098 343440 235060 343496
rect 232037 343438 235060 343440
rect 451444 343496 454007 343498
rect 451444 343440 453946 343496
rect 454002 343440 454007 343496
rect 451444 343438 454007 343440
rect 232037 343435 232103 343438
rect 453941 343435 454007 343438
rect 231945 342138 232011 342141
rect 453941 342138 454007 342141
rect 231945 342136 235060 342138
rect 231945 342080 231950 342136
rect 232006 342080 235060 342136
rect 231945 342078 235060 342080
rect 451444 342136 454007 342138
rect 451444 342080 453946 342136
rect 454002 342080 454007 342136
rect 451444 342078 454007 342080
rect 231945 342075 232011 342078
rect 453941 342075 454007 342078
rect 450854 341396 450860 341460
rect 450924 341458 450930 341460
rect 454033 341458 454099 341461
rect 450924 341456 454099 341458
rect 450924 341400 454038 341456
rect 454094 341400 454099 341456
rect 450924 341398 454099 341400
rect 450924 341396 450930 341398
rect 454033 341395 454099 341398
rect 232037 340778 232103 340781
rect 232037 340776 235060 340778
rect 232037 340720 232042 340776
rect 232098 340720 235060 340776
rect 232037 340718 235060 340720
rect 232037 340715 232103 340718
rect 232221 339962 232287 339965
rect 328494 339962 328500 339964
rect 232221 339960 328500 339962
rect 232221 339904 232226 339960
rect 232282 339904 328500 339960
rect 232221 339902 328500 339904
rect 232221 339899 232287 339902
rect 328494 339900 328500 339902
rect 328564 339900 328570 339964
rect 391790 339900 391796 339964
rect 391860 339962 391866 339964
rect 451038 339962 451044 339964
rect 391860 339902 451044 339962
rect 391860 339900 391866 339902
rect 451038 339900 451044 339902
rect 451108 339900 451114 339964
rect 232497 339826 232563 339829
rect 237414 339826 237420 339828
rect 232497 339824 237420 339826
rect 232497 339768 232502 339824
rect 232558 339768 237420 339824
rect 232497 339766 237420 339768
rect 232497 339763 232563 339766
rect 237414 339764 237420 339766
rect 237484 339764 237490 339828
rect 450118 339764 450124 339828
rect 450188 339826 450194 339828
rect 451230 339826 451290 340748
rect 450188 339766 451290 339826
rect 450188 339764 450194 339766
rect 447726 339628 447732 339692
rect 447796 339690 447802 339692
rect 458357 339690 458423 339693
rect 447796 339688 458423 339690
rect 447796 339632 458362 339688
rect 458418 339632 458423 339688
rect 447796 339630 458423 339632
rect 447796 339628 447802 339630
rect 458357 339627 458423 339630
rect 232037 339418 232103 339421
rect 232037 339416 235060 339418
rect 232037 339360 232042 339416
rect 232098 339360 235060 339416
rect 232037 339358 235060 339360
rect 232037 339355 232103 339358
rect 228449 339282 228515 339285
rect 457529 339282 457595 339285
rect 228449 339280 457595 339282
rect 228449 339224 228454 339280
rect 228510 339224 457534 339280
rect 457590 339224 457595 339280
rect 228449 339222 457595 339224
rect 228449 339219 228515 339222
rect 457529 339219 457595 339222
rect 220445 339010 220511 339013
rect 237230 339010 237236 339012
rect 220445 339008 237236 339010
rect 220445 338952 220450 339008
rect 220506 338952 237236 339008
rect 220445 338950 237236 338952
rect 220445 338947 220511 338950
rect 237230 338948 237236 338950
rect 237300 338948 237306 339012
rect 412398 338948 412404 339012
rect 412468 339010 412474 339012
rect 461669 339010 461735 339013
rect 412468 339008 461735 339010
rect 412468 338952 461674 339008
rect 461730 338952 461735 339008
rect 412468 338950 461735 338952
rect 412468 338948 412474 338950
rect 461669 338947 461735 338950
rect 229921 338874 229987 338877
rect 262806 338874 262812 338876
rect 229921 338872 262812 338874
rect 229921 338816 229926 338872
rect 229982 338816 262812 338872
rect 229921 338814 262812 338816
rect 229921 338811 229987 338814
rect 262806 338812 262812 338814
rect 262876 338812 262882 338876
rect 398966 338812 398972 338876
rect 399036 338874 399042 338876
rect 457069 338874 457135 338877
rect 399036 338872 457135 338874
rect 399036 338816 457074 338872
rect 457130 338816 457135 338872
rect 399036 338814 457135 338816
rect 399036 338812 399042 338814
rect 457069 338811 457135 338814
rect 226793 338738 226859 338741
rect 269246 338738 269252 338740
rect 226793 338736 269252 338738
rect 226793 338680 226798 338736
rect 226854 338680 269252 338736
rect 226793 338678 269252 338680
rect 226793 338675 226859 338678
rect 269246 338676 269252 338678
rect 269316 338676 269322 338740
rect 379646 338676 379652 338740
rect 379716 338738 379722 338740
rect 460381 338738 460447 338741
rect 379716 338736 460447 338738
rect 379716 338680 460386 338736
rect 460442 338680 460447 338736
rect 379716 338678 460447 338680
rect 379716 338676 379722 338678
rect 460381 338675 460447 338678
rect 225689 338602 225755 338605
rect 458817 338602 458883 338605
rect 225689 338600 458883 338602
rect 225689 338544 225694 338600
rect 225750 338544 458822 338600
rect 458878 338544 458883 338600
rect 225689 338542 458883 338544
rect 225689 338539 225755 338542
rect 458817 338539 458883 338542
rect 583520 338452 584960 338692
rect 453573 338330 453639 338333
rect 450494 338328 453639 338330
rect 450494 338272 453578 338328
rect 453634 338272 453639 338328
rect 450494 338270 453639 338272
rect 234245 338194 234311 338197
rect 240501 338194 240567 338197
rect 234245 338192 240567 338194
rect 234245 338136 234250 338192
rect 234306 338136 240506 338192
rect 240562 338136 240567 338192
rect 234245 338134 240567 338136
rect 234245 338131 234311 338134
rect 240501 338131 240567 338134
rect 262806 338132 262812 338196
rect 262876 338194 262882 338196
rect 267733 338194 267799 338197
rect 262876 338192 267799 338194
rect 262876 338136 267738 338192
rect 267794 338136 267799 338192
rect 262876 338134 267799 338136
rect 262876 338132 262882 338134
rect 267733 338131 267799 338134
rect 269246 338132 269252 338196
rect 269316 338194 269322 338196
rect 270769 338194 270835 338197
rect 269316 338192 270835 338194
rect 269316 338136 270774 338192
rect 270830 338136 270835 338192
rect 269316 338134 270835 338136
rect 269316 338132 269322 338134
rect 270769 338131 270835 338134
rect 379513 338194 379579 338197
rect 398925 338196 398991 338197
rect 412357 338196 412423 338197
rect 379646 338194 379652 338196
rect 379513 338192 379652 338194
rect 379513 338136 379518 338192
rect 379574 338136 379652 338192
rect 379513 338134 379652 338136
rect 379513 338131 379579 338134
rect 379646 338132 379652 338134
rect 379716 338132 379722 338196
rect 398925 338194 398972 338196
rect 398880 338192 398972 338194
rect 398880 338136 398930 338192
rect 398880 338134 398972 338136
rect 398925 338132 398972 338134
rect 399036 338132 399042 338196
rect 412357 338194 412404 338196
rect 412312 338192 412404 338194
rect 412312 338136 412362 338192
rect 412312 338134 412404 338136
rect 412357 338132 412404 338134
rect 412468 338132 412474 338196
rect 450353 338194 450419 338197
rect 450494 338194 450554 338270
rect 453573 338267 453639 338270
rect 450353 338192 450554 338194
rect 450353 338136 450358 338192
rect 450414 338136 450554 338192
rect 450353 338134 450554 338136
rect 398925 338131 398991 338132
rect 412357 338131 412423 338132
rect 450353 338131 450419 338134
rect 237230 337860 237236 337924
rect 237300 337922 237306 337924
rect 237373 337922 237439 337925
rect 237300 337920 237439 337922
rect 237300 337864 237378 337920
rect 237434 337864 237439 337920
rect 237300 337862 237439 337864
rect 237300 337860 237306 337862
rect 237373 337859 237439 337862
rect 226190 337588 226196 337652
rect 226260 337650 226266 337652
rect 238753 337650 238819 337653
rect 226260 337648 238819 337650
rect 226260 337592 238758 337648
rect 238814 337592 238819 337648
rect 226260 337590 238819 337592
rect 226260 337588 226266 337590
rect 238753 337587 238819 337590
rect 449893 337650 449959 337653
rect 450862 337650 450922 338028
rect 449893 337648 450922 337650
rect 449893 337592 449898 337648
rect 449954 337592 450922 337648
rect 449893 337590 450922 337592
rect 449893 337587 449959 337590
rect 237414 337452 237420 337516
rect 237484 337514 237490 337516
rect 318793 337514 318859 337517
rect 237484 337512 318859 337514
rect 237484 337456 318798 337512
rect 318854 337456 318859 337512
rect 237484 337454 318859 337456
rect 237484 337452 237490 337454
rect 318793 337451 318859 337454
rect 358813 337514 358879 337517
rect 463969 337514 464035 337517
rect 358813 337512 464035 337514
rect 358813 337456 358818 337512
rect 358874 337456 463974 337512
rect 464030 337456 464035 337512
rect 358813 337454 464035 337456
rect 358813 337451 358879 337454
rect 463969 337451 464035 337454
rect 232814 337316 232820 337380
rect 232884 337378 232890 337380
rect 367737 337378 367803 337381
rect 232884 337376 367803 337378
rect 232884 337320 367742 337376
rect 367798 337320 367803 337376
rect 232884 337318 367803 337320
rect 232884 337316 232890 337318
rect 367737 337315 367803 337318
rect 235390 336636 235396 336700
rect 235460 336698 235466 336700
rect 316033 336698 316099 336701
rect 235460 336696 316099 336698
rect 235460 336640 316038 336696
rect 316094 336640 316099 336696
rect 235460 336638 316099 336640
rect 235460 336636 235466 336638
rect 316033 336635 316099 336638
rect 302233 336562 302299 336565
rect 461158 336562 461164 336564
rect 302233 336560 461164 336562
rect 302233 336504 302238 336560
rect 302294 336504 461164 336560
rect 302233 336502 461164 336504
rect 302233 336499 302299 336502
rect 461158 336500 461164 336502
rect 461228 336500 461234 336564
rect 186313 336426 186379 336429
rect 465441 336426 465507 336429
rect 186313 336424 465507 336426
rect 186313 336368 186318 336424
rect 186374 336368 465446 336424
rect 465502 336368 465507 336424
rect 186313 336366 465507 336368
rect 186313 336363 186379 336366
rect 465441 336363 465507 336366
rect 182173 336290 182239 336293
rect 461342 336290 461348 336292
rect 182173 336288 461348 336290
rect 182173 336232 182178 336288
rect 182234 336232 461348 336288
rect 182173 336230 461348 336232
rect 182173 336227 182239 336230
rect 461342 336228 461348 336230
rect 461412 336228 461418 336292
rect 171133 336154 171199 336157
rect 459502 336154 459508 336156
rect 171133 336152 459508 336154
rect 171133 336096 171138 336152
rect 171194 336096 459508 336152
rect 171133 336094 459508 336096
rect 171133 336091 171199 336094
rect 459502 336092 459508 336094
rect 459572 336092 459578 336156
rect 146293 336018 146359 336021
rect 460105 336018 460171 336021
rect 146293 336016 460171 336018
rect 146293 335960 146298 336016
rect 146354 335960 460110 336016
rect 460166 335960 460171 336016
rect 146293 335958 460171 335960
rect 146293 335955 146359 335958
rect 460105 335955 460171 335958
rect 157333 334658 157399 334661
rect 462262 334658 462268 334660
rect 157333 334656 462268 334658
rect 157333 334600 157338 334656
rect 157394 334600 462268 334656
rect 157333 334598 462268 334600
rect 157333 334595 157399 334598
rect 462262 334596 462268 334598
rect 462332 334596 462338 334660
rect 441613 334114 441679 334117
rect 450118 334114 450124 334116
rect 441613 334112 450124 334114
rect 441613 334056 441618 334112
rect 441674 334056 450124 334112
rect 441613 334054 450124 334056
rect 441613 334051 441679 334054
rect 450118 334052 450124 334054
rect 450188 334052 450194 334116
rect 124213 333570 124279 333573
rect 463734 333570 463740 333572
rect 124213 333568 463740 333570
rect 124213 333512 124218 333568
rect 124274 333512 463740 333568
rect 124213 333510 463740 333512
rect 124213 333507 124279 333510
rect 463734 333508 463740 333510
rect 463804 333508 463810 333572
rect 63493 333434 63559 333437
rect 458909 333434 458975 333437
rect 63493 333432 458975 333434
rect 63493 333376 63498 333432
rect 63554 333376 458914 333432
rect 458970 333376 458975 333432
rect 63493 333374 458975 333376
rect 63493 333371 63559 333374
rect 458909 333371 458975 333374
rect 19333 333298 19399 333301
rect 465533 333298 465599 333301
rect 19333 333296 465599 333298
rect 19333 333240 19338 333296
rect 19394 333240 465538 333296
rect 465594 333240 465599 333296
rect 19333 333238 465599 333240
rect 19333 333235 19399 333238
rect 465533 333235 465599 333238
rect 227110 333100 227116 333164
rect 227180 333162 227186 333164
rect 230473 333162 230539 333165
rect 227180 333160 230539 333162
rect 227180 333104 230478 333160
rect 230534 333104 230539 333160
rect 227180 333102 230539 333104
rect 227180 333100 227186 333102
rect 230473 333099 230539 333102
rect -960 332196 480 332436
rect 233182 331740 233188 331804
rect 233252 331802 233258 331804
rect 505093 331802 505159 331805
rect 233252 331800 505159 331802
rect 233252 331744 505098 331800
rect 505154 331744 505159 331800
rect 233252 331742 505159 331744
rect 233252 331740 233258 331742
rect 505093 331739 505159 331742
rect 229870 330380 229876 330444
rect 229940 330442 229946 330444
rect 578233 330442 578299 330445
rect 229940 330440 578299 330442
rect 229940 330384 578238 330440
rect 578294 330384 578299 330440
rect 229940 330382 578299 330384
rect 229940 330380 229946 330382
rect 578233 330379 578299 330382
rect 233366 329156 233372 329220
rect 233436 329218 233442 329220
rect 507853 329218 507919 329221
rect 233436 329216 507919 329218
rect 233436 329160 507858 329216
rect 507914 329160 507919 329216
rect 233436 329158 507919 329160
rect 233436 329156 233442 329158
rect 507853 329155 507919 329158
rect 230054 329020 230060 329084
rect 230124 329082 230130 329084
rect 517513 329082 517579 329085
rect 230124 329080 517579 329082
rect 230124 329024 517518 329080
rect 517574 329024 517579 329080
rect 230124 329022 517579 329024
rect 230124 329020 230130 329022
rect 517513 329019 517579 329022
rect 235022 327796 235028 327860
rect 235092 327858 235098 327860
rect 266353 327858 266419 327861
rect 235092 327856 266419 327858
rect 235092 327800 266358 327856
rect 266414 327800 266419 327856
rect 235092 327798 266419 327800
rect 235092 327796 235098 327798
rect 266353 327795 266419 327798
rect 5533 327722 5599 327725
rect 457110 327722 457116 327724
rect 5533 327720 457116 327722
rect 5533 327664 5538 327720
rect 5594 327664 457116 327720
rect 5533 327662 457116 327664
rect 5533 327659 5599 327662
rect 457110 327660 457116 327662
rect 457180 327660 457186 327724
rect 228766 326300 228772 326364
rect 228836 326362 228842 326364
rect 390553 326362 390619 326365
rect 228836 326360 390619 326362
rect 228836 326304 390558 326360
rect 390614 326304 390619 326360
rect 228836 326302 390619 326304
rect 228836 326300 228842 326302
rect 390553 326299 390619 326302
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 212533 323778 212599 323781
rect 455638 323778 455644 323780
rect 212533 323776 455644 323778
rect 212533 323720 212538 323776
rect 212594 323720 455644 323776
rect 212533 323718 455644 323720
rect 212533 323715 212599 323718
rect 455638 323716 455644 323718
rect 455708 323716 455714 323780
rect 110413 323642 110479 323645
rect 451406 323642 451412 323644
rect 110413 323640 451412 323642
rect 110413 323584 110418 323640
rect 110474 323584 451412 323640
rect 110413 323582 451412 323584
rect 110413 323579 110479 323582
rect 451406 323580 451412 323582
rect 451476 323580 451482 323644
rect 35893 322146 35959 322149
rect 458766 322146 458772 322148
rect 35893 322144 458772 322146
rect 35893 322088 35898 322144
rect 35954 322088 458772 322144
rect 35893 322086 458772 322088
rect 35893 322083 35959 322086
rect 458766 322084 458772 322086
rect 458836 322084 458842 322148
rect 75913 320922 75979 320925
rect 457294 320922 457300 320924
rect 75913 320920 457300 320922
rect 75913 320864 75918 320920
rect 75974 320864 457300 320920
rect 75913 320862 457300 320864
rect 75913 320859 75979 320862
rect 457294 320860 457300 320862
rect 457364 320860 457370 320924
rect 13 320786 79 320789
rect 450302 320786 450308 320788
rect 13 320784 450308 320786
rect 13 320728 18 320784
rect 74 320728 450308 320784
rect 13 320726 450308 320728
rect 13 320723 79 320726
rect 450302 320724 450308 320726
rect 450372 320724 450378 320788
rect -960 319290 480 319380
rect 3509 319290 3575 319293
rect -960 319288 3575 319290
rect -960 319232 3514 319288
rect 3570 319232 3575 319288
rect -960 319230 3575 319232
rect -960 319140 480 319230
rect 3509 319227 3575 319230
rect 232446 318140 232452 318204
rect 232516 318202 232522 318204
rect 552013 318202 552079 318205
rect 232516 318200 552079 318202
rect 232516 318144 552018 318200
rect 552074 318144 552079 318200
rect 232516 318142 552079 318144
rect 232516 318140 232522 318142
rect 552013 318139 552079 318142
rect 235206 318004 235212 318068
rect 235276 318066 235282 318068
rect 580993 318066 581059 318069
rect 235276 318064 581059 318066
rect 235276 318008 580998 318064
rect 581054 318008 581059 318064
rect 235276 318006 581059 318008
rect 235276 318004 235282 318006
rect 580993 318003 581059 318006
rect 228582 316916 228588 316980
rect 228652 316978 228658 316980
rect 382365 316978 382431 316981
rect 228652 316976 382431 316978
rect 228652 316920 382370 316976
rect 382426 316920 382431 316976
rect 228652 316918 382431 316920
rect 228652 316916 228658 316918
rect 382365 316915 382431 316918
rect 232630 316780 232636 316844
rect 232700 316842 232706 316844
rect 523125 316842 523191 316845
rect 232700 316840 523191 316842
rect 232700 316784 523130 316840
rect 523186 316784 523191 316840
rect 232700 316782 523191 316784
rect 232700 316780 232706 316782
rect 523125 316779 523191 316782
rect 44265 316706 44331 316709
rect 456006 316706 456012 316708
rect 44265 316704 456012 316706
rect 44265 316648 44270 316704
rect 44326 316648 456012 316704
rect 44265 316646 456012 316648
rect 44265 316643 44331 316646
rect 456006 316644 456012 316646
rect 456076 316644 456082 316708
rect 71773 315346 71839 315349
rect 456926 315346 456932 315348
rect 71773 315344 456932 315346
rect 71773 315288 71778 315344
rect 71834 315288 456932 315344
rect 71773 315286 456932 315288
rect 71773 315283 71839 315286
rect 456926 315284 456932 315286
rect 456996 315284 457002 315348
rect 60825 314122 60891 314125
rect 452878 314122 452884 314124
rect 60825 314120 452884 314122
rect 60825 314064 60830 314120
rect 60886 314064 452884 314120
rect 60825 314062 452884 314064
rect 60825 314059 60891 314062
rect 452878 314060 452884 314062
rect 452948 314060 452954 314124
rect 41413 313986 41479 313989
rect 458582 313986 458588 313988
rect 41413 313984 458588 313986
rect 41413 313928 41418 313984
rect 41474 313928 458588 313984
rect 41413 313926 458588 313928
rect 41413 313923 41479 313926
rect 458582 313924 458588 313926
rect 458652 313924 458658 313988
rect 22093 312490 22159 312493
rect 453246 312490 453252 312492
rect 22093 312488 453252 312490
rect 22093 312432 22098 312488
rect 22154 312432 453252 312488
rect 22093 312430 453252 312432
rect 22093 312427 22159 312430
rect 453246 312428 453252 312430
rect 453316 312428 453322 312492
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 97993 311130 98059 311133
rect 454534 311130 454540 311132
rect 97993 311128 454540 311130
rect 97993 311072 97998 311128
rect 98054 311072 454540 311128
rect 97993 311070 454540 311072
rect 97993 311067 98059 311070
rect 454534 311068 454540 311070
rect 454604 311068 454610 311132
rect 56593 309770 56659 309773
rect 458398 309770 458404 309772
rect 56593 309768 458404 309770
rect 56593 309712 56598 309768
rect 56654 309712 458404 309768
rect 56593 309710 458404 309712
rect 56593 309707 56659 309710
rect 458398 309708 458404 309710
rect 458468 309708 458474 309772
rect 180793 308410 180859 308413
rect 453062 308410 453068 308412
rect 180793 308408 453068 308410
rect 180793 308352 180798 308408
rect 180854 308352 453068 308408
rect 180793 308350 453068 308352
rect 180793 308347 180859 308350
rect 453062 308348 453068 308350
rect 453132 308348 453138 308412
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 230238 304132 230244 304196
rect 230308 304194 230314 304196
rect 445753 304194 445819 304197
rect 230308 304192 445819 304194
rect 230308 304136 445758 304192
rect 445814 304136 445819 304192
rect 230308 304134 445819 304136
rect 230308 304132 230314 304134
rect 445753 304131 445819 304134
rect 135253 301474 135319 301477
rect 454350 301474 454356 301476
rect 135253 301472 454356 301474
rect 135253 301416 135258 301472
rect 135314 301416 454356 301472
rect 135253 301414 454356 301416
rect 135253 301411 135319 301414
rect 454350 301412 454356 301414
rect 454420 301412 454426 301476
rect 231158 300052 231164 300116
rect 231228 300114 231234 300116
rect 456793 300114 456859 300117
rect 231228 300112 456859 300114
rect 231228 300056 456798 300112
rect 456854 300056 456859 300112
rect 231228 300054 456859 300056
rect 231228 300052 231234 300054
rect 456793 300051 456859 300054
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 118785 296034 118851 296037
rect 455822 296034 455828 296036
rect 118785 296032 455828 296034
rect 118785 295976 118790 296032
rect 118846 295976 455828 296032
rect 118785 295974 455828 295976
rect 118785 295971 118851 295974
rect 455822 295972 455828 295974
rect 455892 295972 455898 296036
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 232998 293116 233004 293180
rect 233068 293178 233074 293180
rect 447777 293178 447843 293181
rect 233068 293176 447843 293178
rect 233068 293120 447782 293176
rect 447838 293120 447843 293176
rect 233068 293118 447843 293120
rect 233068 293116 233074 293118
rect 447777 293115 447843 293118
rect 583520 285276 584960 285516
rect 93853 283522 93919 283525
rect 458214 283522 458220 283524
rect 93853 283520 458220 283522
rect 93853 283464 93858 283520
rect 93914 283464 458220 283520
rect 93853 283462 458220 283464
rect 93853 283459 93919 283462
rect 458214 283460 458220 283462
rect 458284 283460 458290 283524
rect -960 279972 480 280212
rect 227294 279380 227300 279444
rect 227364 279442 227370 279444
rect 581085 279442 581151 279445
rect 227364 279440 581151 279442
rect 227364 279384 581090 279440
rect 581146 279384 581151 279440
rect 227364 279382 581151 279384
rect 227364 279380 227370 279382
rect 581085 279379 581151 279382
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 227478 261428 227484 261492
rect 227548 261490 227554 261492
rect 456885 261490 456951 261493
rect 227548 261488 456951 261490
rect 227548 261432 456890 261488
rect 456946 261432 456951 261488
rect 227548 261430 456951 261432
rect 227548 261428 227554 261430
rect 456885 261427 456951 261430
rect 580625 258906 580691 258909
rect 583520 258906 584960 258996
rect 580625 258904 584960 258906
rect 580625 258848 580630 258904
rect 580686 258848 584960 258904
rect 580625 258846 584960 258848
rect 580625 258843 580691 258846
rect 233550 258708 233556 258772
rect 233620 258770 233626 258772
rect 580441 258770 580507 258773
rect 233620 258768 580507 258770
rect 233620 258712 580446 258768
rect 580502 258712 580507 258768
rect 583520 258756 584960 258846
rect 233620 258710 580507 258712
rect 233620 258708 233626 258710
rect 580441 258707 580507 258710
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 64873 251834 64939 251837
rect 456742 251834 456748 251836
rect 64873 251832 456748 251834
rect 64873 251776 64878 251832
rect 64934 251776 456748 251832
rect 64873 251774 456748 251776
rect 64873 251771 64939 251774
rect 456742 251772 456748 251774
rect 456812 251772 456818 251836
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 580349 232386 580415 232389
rect 583520 232386 584960 232476
rect 580349 232384 584960 232386
rect 580349 232328 580354 232384
rect 580410 232328 584960 232384
rect 580349 232326 584960 232328
rect 580349 232323 580415 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579981 205730 580047 205733
rect 583520 205730 584960 205820
rect 579981 205728 584960 205730
rect 579981 205672 579986 205728
rect 580042 205672 584960 205728
rect 579981 205670 584960 205672
rect 579981 205667 580047 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 231342 170308 231348 170372
rect 231412 170370 231418 170372
rect 521653 170370 521719 170373
rect 231412 170368 521719 170370
rect 231412 170312 521658 170368
rect 521714 170312 521719 170368
rect 231412 170310 521719 170312
rect 231412 170308 231418 170310
rect 521653 170307 521719 170310
rect 2865 166290 2931 166293
rect 454166 166290 454172 166292
rect 2865 166288 454172 166290
rect 2865 166232 2870 166288
rect 2926 166232 454172 166288
rect 2865 166230 454172 166232
rect 2865 166227 2931 166230
rect 454166 166228 454172 166230
rect 454236 166228 454242 166292
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 225638 136778 225644 136780
rect -960 136718 225644 136778
rect -960 136628 480 136718
rect 225638 136716 225644 136718
rect 225708 136716 225714 136780
rect 580257 126034 580323 126037
rect 583520 126034 584960 126124
rect 580257 126032 584960 126034
rect 580257 125976 580262 126032
rect 580318 125976 584960 126032
rect 580257 125974 584960 125976
rect 580257 125971 580323 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 154573 112434 154639 112437
rect 455454 112434 455460 112436
rect 154573 112432 455460 112434
rect 154573 112376 154578 112432
rect 154634 112376 455460 112432
rect 154573 112374 455460 112376
rect 154573 112371 154639 112374
rect 455454 112372 455460 112374
rect 455524 112372 455530 112436
rect 233734 111828 233740 111892
rect 233804 111890 233810 111892
rect 583526 111890 583586 112646
rect 233804 111830 583586 111890
rect 233804 111828 233810 111830
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580441 59666 580507 59669
rect 583520 59666 584960 59756
rect 580441 59664 584960 59666
rect 580441 59608 580446 59664
rect 580502 59608 584960 59664
rect 580441 59606 584960 59608
rect 580441 59603 580507 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect -960 58518 674 58578
rect -960 58442 480 58518
rect 614 58442 674 58518
rect -960 58428 674 58442
rect 246 58382 674 58428
rect 246 58034 306 58382
rect 228214 58034 228220 58036
rect 246 57974 228220 58034
rect 228214 57972 228220 57974
rect 228284 57972 228290 58036
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 231710 37844 231716 37908
rect 231780 37906 231786 37908
rect 476113 37906 476179 37909
rect 231780 37904 476179 37906
rect 231780 37848 476118 37904
rect 476174 37848 476179 37904
rect 231780 37846 476179 37848
rect 231780 37844 231786 37846
rect 476113 37843 476179 37846
rect 231526 36484 231532 36548
rect 231596 36546 231602 36548
rect 465257 36546 465323 36549
rect 231596 36544 465323 36546
rect 231596 36488 465262 36544
rect 465318 36488 465323 36544
rect 231596 36486 465323 36488
rect 231596 36484 231602 36486
rect 465257 36483 465323 36486
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 93945 15874 94011 15877
rect 452694 15874 452700 15876
rect 93945 15872 452700 15874
rect 93945 15816 93950 15872
rect 94006 15816 452700 15872
rect 93945 15814 452700 15816
rect 93945 15811 94011 15814
rect 452694 15812 452700 15814
rect 452764 15812 452770 15876
rect 184933 11658 184999 11661
rect 454166 11658 454172 11660
rect 184933 11656 454172 11658
rect 184933 11600 184938 11656
rect 184994 11600 454172 11656
rect 184933 11598 454172 11600
rect 184933 11595 184999 11598
rect 454166 11596 454172 11598
rect 454236 11596 454242 11660
rect 223297 6626 223363 6629
rect 310237 6626 310303 6629
rect 223297 6624 310303 6626
rect -960 6490 480 6580
rect 223297 6568 223302 6624
rect 223358 6568 310242 6624
rect 310298 6568 310303 6624
rect 223297 6566 310303 6568
rect 223297 6563 223363 6566
rect 310237 6563 310303 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 213821 6490 213887 6493
rect 356329 6490 356395 6493
rect 213821 6488 356395 6490
rect 213821 6432 213826 6488
rect 213882 6432 356334 6488
rect 356390 6432 356395 6488
rect 213821 6430 356395 6432
rect 213821 6427 213887 6430
rect 356329 6427 356395 6430
rect 365805 6490 365871 6493
rect 450486 6490 450492 6492
rect 365805 6488 450492 6490
rect 365805 6432 365810 6488
rect 365866 6432 450492 6488
rect 365805 6430 450492 6432
rect 365805 6427 365871 6430
rect 450486 6428 450492 6430
rect 450556 6428 450562 6492
rect 583520 6476 584960 6566
rect 230105 6354 230171 6357
rect 559741 6354 559807 6357
rect 230105 6352 559807 6354
rect 230105 6296 230110 6352
rect 230166 6296 559746 6352
rect 559802 6296 559807 6352
rect 230105 6294 559807 6296
rect 230105 6291 230171 6294
rect 559741 6291 559807 6294
rect 224401 6218 224467 6221
rect 553761 6218 553827 6221
rect 224401 6216 553827 6218
rect 224401 6160 224406 6216
rect 224462 6160 553766 6216
rect 553822 6160 553827 6216
rect 224401 6158 553827 6160
rect 224401 6155 224467 6158
rect 553761 6155 553827 6158
rect 179045 4042 179111 4045
rect 225454 4042 225460 4044
rect 179045 4040 225460 4042
rect 179045 3984 179050 4040
rect 179106 3984 225460 4040
rect 179045 3982 225460 3984
rect 179045 3979 179111 3982
rect 225454 3980 225460 3982
rect 225524 3980 225530 4044
rect 228950 3980 228956 4044
rect 229020 4042 229026 4044
rect 337469 4042 337535 4045
rect 229020 4040 337535 4042
rect 229020 3984 337474 4040
rect 337530 3984 337535 4040
rect 229020 3982 337535 3984
rect 229020 3980 229026 3982
rect 337469 3979 337535 3982
rect 351637 4042 351703 4045
rect 447726 4042 447732 4044
rect 351637 4040 447732 4042
rect 351637 3984 351642 4040
rect 351698 3984 447732 4040
rect 351637 3982 447732 3984
rect 351637 3979 351703 3982
rect 447726 3980 447732 3982
rect 447796 3980 447802 4044
rect 138841 3906 138907 3909
rect 229686 3906 229692 3908
rect 138841 3904 229692 3906
rect 138841 3848 138846 3904
rect 138902 3848 229692 3904
rect 138841 3846 229692 3848
rect 138841 3843 138907 3846
rect 229686 3844 229692 3846
rect 229756 3844 229762 3908
rect 327993 3906 328059 3909
rect 451958 3906 451964 3908
rect 327993 3904 451964 3906
rect 327993 3848 327998 3904
rect 328054 3848 451964 3904
rect 327993 3846 451964 3848
rect 327993 3843 328059 3846
rect 451958 3844 451964 3846
rect 452028 3844 452034 3908
rect 224769 3770 224835 3773
rect 530117 3770 530183 3773
rect 224769 3768 530183 3770
rect 224769 3712 224774 3768
rect 224830 3712 530122 3768
rect 530178 3712 530183 3768
rect 224769 3710 530183 3712
rect 224769 3707 224835 3710
rect 530117 3707 530183 3710
rect 39573 3634 39639 3637
rect 364425 3634 364491 3637
rect 39573 3632 364491 3634
rect 39573 3576 39578 3632
rect 39634 3576 364430 3632
rect 364486 3576 364491 3632
rect 39573 3574 364491 3576
rect 39573 3571 39639 3574
rect 364425 3571 364491 3574
rect 436737 3634 436803 3637
rect 465901 3634 465967 3637
rect 436737 3632 465967 3634
rect 436737 3576 436742 3632
rect 436798 3576 465906 3632
rect 465962 3576 465967 3632
rect 436737 3574 465967 3576
rect 436737 3571 436803 3574
rect 465901 3571 465967 3574
rect 32397 3498 32463 3501
rect 363045 3498 363111 3501
rect 391841 3500 391907 3501
rect 32397 3496 363111 3498
rect 32397 3440 32402 3496
rect 32458 3440 363050 3496
rect 363106 3440 363111 3496
rect 32397 3438 363111 3440
rect 32397 3435 32463 3438
rect 363045 3435 363111 3438
rect 391790 3436 391796 3500
rect 391860 3498 391907 3500
rect 391860 3496 391952 3498
rect 391902 3440 391952 3496
rect 391860 3438 391952 3440
rect 391860 3436 391907 3438
rect 460054 3436 460060 3500
rect 460124 3498 460130 3500
rect 568021 3498 568087 3501
rect 460124 3496 568087 3498
rect 460124 3440 568026 3496
rect 568082 3440 568087 3496
rect 460124 3438 568087 3440
rect 460124 3436 460130 3438
rect 391841 3435 391907 3436
rect 568021 3435 568087 3438
rect 20621 3362 20687 3365
rect 381537 3362 381603 3365
rect 20621 3360 381603 3362
rect 20621 3304 20626 3360
rect 20682 3304 381542 3360
rect 381598 3304 381603 3360
rect 20621 3302 381603 3304
rect 20621 3299 20687 3302
rect 381537 3299 381603 3302
rect 460238 3300 460244 3364
rect 460308 3362 460314 3364
rect 583385 3362 583451 3365
rect 460308 3360 583451 3362
rect 460308 3304 583390 3360
rect 583446 3304 583451 3360
rect 460308 3302 583451 3304
rect 460308 3300 460314 3302
rect 583385 3299 583451 3302
rect 328494 3164 328500 3228
rect 328564 3226 328570 3228
rect 329189 3226 329255 3229
rect 328564 3224 329255 3226
rect 328564 3168 329194 3224
rect 329250 3168 329255 3224
rect 328564 3166 329255 3168
rect 328564 3164 328570 3166
rect 329189 3163 329255 3166
rect 437933 3226 437999 3229
rect 463785 3226 463851 3229
rect 437933 3224 463851 3226
rect 437933 3168 437938 3224
rect 437994 3168 463790 3224
rect 463846 3168 463851 3224
rect 437933 3166 463851 3168
rect 437933 3163 437999 3166
rect 463785 3163 463851 3166
<< via3 >>
rect 460980 632028 461044 632092
rect 225644 560492 225708 560556
rect 227116 560356 227180 560420
rect 226196 559812 226260 559876
rect 461164 558996 461228 559060
rect 229692 558044 229756 558108
rect 228220 557908 228284 557972
rect 460060 557772 460124 557836
rect 228956 556820 229020 556884
rect 451044 556820 451108 556884
rect 235764 556684 235828 556748
rect 460244 556548 460308 556612
rect 225460 556412 225524 556476
rect 264652 555928 264716 555932
rect 264652 555872 264656 555928
rect 264656 555872 264712 555928
rect 264712 555872 264716 555928
rect 264652 555868 264716 555872
rect 352236 555928 352300 555932
rect 352236 555872 352240 555928
rect 352240 555872 352296 555928
rect 352296 555872 352300 555928
rect 352236 555868 352300 555872
rect 264652 555188 264716 555252
rect 352236 554780 352300 554844
rect 235764 554508 235828 554572
rect 458404 552876 458468 552940
rect 455644 551516 455708 551580
rect 231164 550156 231228 550220
rect 458588 548796 458652 548860
rect 227300 542404 227364 542468
rect 452884 539276 452948 539340
rect 231348 535876 231412 535940
rect 227484 531388 227548 531452
rect 458220 529076 458284 529140
rect 230244 527716 230308 527780
rect 233372 523636 233436 523700
rect 456748 523636 456812 523700
rect 228772 517516 228836 517580
rect 230060 513436 230124 513500
rect 231716 512076 231780 512140
rect 463740 510580 463804 510644
rect 461348 506500 461412 506564
rect 456932 505276 456996 505340
rect 233740 503916 233804 503980
rect 458772 501196 458836 501260
rect 231532 497796 231596 497860
rect 454172 497116 454236 497180
rect 451412 493716 451476 493780
rect 228588 491268 228652 491332
rect 459508 484196 459572 484260
rect 233556 469916 233620 469980
rect 233004 467196 233068 467260
rect 455460 461756 455524 461820
rect 454356 448836 454420 448900
rect 233188 447476 233252 447540
rect 454172 446116 454236 446180
rect 457116 443396 457180 443460
rect 462268 441628 462332 441692
rect 232820 437276 232884 437340
rect 457300 433196 457364 433260
rect 235028 427756 235092 427820
rect 454540 422316 454604 422380
rect 456012 415516 456076 415580
rect 229876 414836 229940 414900
rect 455828 412116 455892 412180
rect 452700 410756 452764 410820
rect 451964 409940 452028 410004
rect 232636 406676 232700 406740
rect 450860 403956 450924 404020
rect 453068 398516 453132 398580
rect 232452 388316 232516 388380
rect 235212 386956 235276 387020
rect 460980 360164 461044 360228
rect 235396 358396 235460 358460
rect 453252 351596 453316 351660
rect 450860 341396 450924 341460
rect 328500 339900 328564 339964
rect 391796 339900 391860 339964
rect 451044 339900 451108 339964
rect 237420 339764 237484 339828
rect 450124 339764 450188 339828
rect 447732 339628 447796 339692
rect 237236 338948 237300 339012
rect 412404 338948 412468 339012
rect 262812 338812 262876 338876
rect 398972 338812 399036 338876
rect 269252 338676 269316 338740
rect 379652 338676 379716 338740
rect 262812 338132 262876 338196
rect 269252 338132 269316 338196
rect 379652 338132 379716 338196
rect 398972 338192 399036 338196
rect 398972 338136 398986 338192
rect 398986 338136 399036 338192
rect 398972 338132 399036 338136
rect 412404 338192 412468 338196
rect 412404 338136 412418 338192
rect 412418 338136 412468 338192
rect 412404 338132 412468 338136
rect 237236 337860 237300 337924
rect 226196 337588 226260 337652
rect 237420 337452 237484 337516
rect 232820 337316 232884 337380
rect 235396 336636 235460 336700
rect 461164 336500 461228 336564
rect 461348 336228 461412 336292
rect 459508 336092 459572 336156
rect 462268 334596 462332 334660
rect 450124 334052 450188 334116
rect 463740 333508 463804 333572
rect 227116 333100 227180 333164
rect 233188 331740 233252 331804
rect 229876 330380 229940 330444
rect 233372 329156 233436 329220
rect 230060 329020 230124 329084
rect 235028 327796 235092 327860
rect 457116 327660 457180 327724
rect 228772 326300 228836 326364
rect 455644 323716 455708 323780
rect 451412 323580 451476 323644
rect 458772 322084 458836 322148
rect 457300 320860 457364 320924
rect 450308 320724 450372 320788
rect 232452 318140 232516 318204
rect 235212 318004 235276 318068
rect 228588 316916 228652 316980
rect 232636 316780 232700 316844
rect 456012 316644 456076 316708
rect 456932 315284 456996 315348
rect 452884 314060 452948 314124
rect 458588 313924 458652 313988
rect 453252 312428 453316 312492
rect 454540 311068 454604 311132
rect 458404 309708 458468 309772
rect 453068 308348 453132 308412
rect 230244 304132 230308 304196
rect 454356 301412 454420 301476
rect 231164 300052 231228 300116
rect 455828 295972 455892 296036
rect 233004 293116 233068 293180
rect 458220 283460 458284 283524
rect 227300 279380 227364 279444
rect 227484 261428 227548 261492
rect 233556 258708 233620 258772
rect 456748 251772 456812 251836
rect 231348 170308 231412 170372
rect 454172 166228 454236 166292
rect 225644 136716 225708 136780
rect 455460 112372 455524 112436
rect 233740 111828 233804 111892
rect 228220 57972 228284 58036
rect 231716 37844 231780 37908
rect 231532 36484 231596 36548
rect 452700 15812 452764 15876
rect 454172 11596 454236 11660
rect 450492 6428 450556 6492
rect 225460 3980 225524 4044
rect 228956 3980 229020 4044
rect 447732 3980 447796 4044
rect 229692 3844 229756 3908
rect 451964 3844 452028 3908
rect 391796 3496 391860 3500
rect 391796 3440 391846 3496
rect 391846 3440 391860 3496
rect 391796 3436 391860 3440
rect 460060 3436 460124 3500
rect 460244 3300 460308 3364
rect 328500 3164 328564 3228
<< metal4 >>
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 705798 6134 705830
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -1894 6134 -1862
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 705798 42134 705830
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -1894 42134 -1862
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 705798 78134 705830
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -1894 78134 -1862
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 705798 114134 705830
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -1894 114134 -1862
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 705798 150134 705830
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -1894 150134 -1862
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 705798 186134 705830
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -1894 186134 -1862
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 705798 222134 705830
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 225643 560556 225709 560557
rect 225643 560492 225644 560556
rect 225708 560492 225709 560556
rect 225643 560491 225709 560492
rect 225459 556476 225525 556477
rect 225459 556412 225460 556476
rect 225524 556412 225525 556476
rect 225459 556411 225525 556412
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 225462 4045 225522 556411
rect 225646 136781 225706 560491
rect 227115 560420 227181 560421
rect 227115 560356 227116 560420
rect 227180 560356 227181 560420
rect 227115 560355 227181 560356
rect 226195 559876 226261 559877
rect 226195 559812 226196 559876
rect 226260 559812 226261 559876
rect 226195 559811 226261 559812
rect 226198 337653 226258 559811
rect 226195 337652 226261 337653
rect 226195 337588 226196 337652
rect 226260 337588 226261 337652
rect 226195 337587 226261 337588
rect 227118 333165 227178 560355
rect 229691 558108 229757 558109
rect 229691 558044 229692 558108
rect 229756 558044 229757 558108
rect 229691 558043 229757 558044
rect 228219 557972 228285 557973
rect 228219 557908 228220 557972
rect 228284 557908 228285 557972
rect 228219 557907 228285 557908
rect 227299 542468 227365 542469
rect 227299 542404 227300 542468
rect 227364 542404 227365 542468
rect 227299 542403 227365 542404
rect 227115 333164 227181 333165
rect 227115 333100 227116 333164
rect 227180 333100 227181 333164
rect 227115 333099 227181 333100
rect 227302 279445 227362 542403
rect 227483 531452 227549 531453
rect 227483 531388 227484 531452
rect 227548 531388 227549 531452
rect 227483 531387 227549 531388
rect 227299 279444 227365 279445
rect 227299 279380 227300 279444
rect 227364 279380 227365 279444
rect 227299 279379 227365 279380
rect 227486 261493 227546 531387
rect 227483 261492 227549 261493
rect 227483 261428 227484 261492
rect 227548 261428 227549 261492
rect 227483 261427 227549 261428
rect 225643 136780 225709 136781
rect 225643 136716 225644 136780
rect 225708 136716 225709 136780
rect 225643 136715 225709 136716
rect 228222 58037 228282 557907
rect 228955 556884 229021 556885
rect 228955 556820 228956 556884
rect 229020 556820 229021 556884
rect 228955 556819 229021 556820
rect 228771 517580 228837 517581
rect 228771 517516 228772 517580
rect 228836 517516 228837 517580
rect 228771 517515 228837 517516
rect 228587 491332 228653 491333
rect 228587 491268 228588 491332
rect 228652 491268 228653 491332
rect 228587 491267 228653 491268
rect 228590 316981 228650 491267
rect 228774 326365 228834 517515
rect 228771 326364 228837 326365
rect 228771 326300 228772 326364
rect 228836 326300 228837 326364
rect 228771 326299 228837 326300
rect 228587 316980 228653 316981
rect 228587 316916 228588 316980
rect 228652 316916 228653 316980
rect 228587 316915 228653 316916
rect 228219 58036 228285 58037
rect 228219 57972 228220 58036
rect 228284 57972 228285 58036
rect 228219 57971 228285 57972
rect 228958 4045 229018 556819
rect 225459 4044 225525 4045
rect 225459 3980 225460 4044
rect 225524 3980 225525 4044
rect 225459 3979 225525 3980
rect 228955 4044 229021 4045
rect 228955 3980 228956 4044
rect 229020 3980 229021 4044
rect 228955 3979 229021 3980
rect 229694 3909 229754 558043
rect 235763 556748 235829 556749
rect 235763 556684 235764 556748
rect 235828 556684 235829 556748
rect 235763 556683 235829 556684
rect 235766 554573 235826 556683
rect 235763 554572 235829 554573
rect 235763 554508 235764 554572
rect 235828 554508 235829 554572
rect 235763 554507 235829 554508
rect 231163 550220 231229 550221
rect 231163 550156 231164 550220
rect 231228 550156 231229 550220
rect 231163 550155 231229 550156
rect 230243 527780 230309 527781
rect 230243 527716 230244 527780
rect 230308 527716 230309 527780
rect 230243 527715 230309 527716
rect 230059 513500 230125 513501
rect 230059 513436 230060 513500
rect 230124 513436 230125 513500
rect 230059 513435 230125 513436
rect 229875 414900 229941 414901
rect 229875 414836 229876 414900
rect 229940 414836 229941 414900
rect 229875 414835 229941 414836
rect 229878 330445 229938 414835
rect 229875 330444 229941 330445
rect 229875 330380 229876 330444
rect 229940 330380 229941 330444
rect 229875 330379 229941 330380
rect 230062 329085 230122 513435
rect 230059 329084 230125 329085
rect 230059 329020 230060 329084
rect 230124 329020 230125 329084
rect 230059 329019 230125 329020
rect 230246 304197 230306 527715
rect 230243 304196 230309 304197
rect 230243 304132 230244 304196
rect 230308 304132 230309 304196
rect 230243 304131 230309 304132
rect 231166 300117 231226 550155
rect 253794 547017 254414 578898
rect 257514 705798 258134 705830
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547017 258134 582618
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 264651 555932 264717 555933
rect 264651 555868 264652 555932
rect 264716 555868 264717 555932
rect 264651 555867 264717 555868
rect 264654 555253 264714 555867
rect 264651 555252 264717 555253
rect 264651 555188 264652 555252
rect 264716 555188 264717 555252
rect 264651 555187 264717 555188
rect 289794 547017 290414 578898
rect 293514 705798 294134 705830
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547017 294134 582618
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 547017 326414 578898
rect 329514 705798 330134 705830
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547017 330134 582618
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 352235 555932 352301 555933
rect 352235 555868 352236 555932
rect 352300 555868 352301 555932
rect 352235 555867 352301 555868
rect 352238 554845 352298 555867
rect 352235 554844 352301 554845
rect 352235 554780 352236 554844
rect 352300 554780 352301 554844
rect 352235 554779 352301 554780
rect 361794 547017 362414 578898
rect 365514 705798 366134 705830
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547017 366134 582618
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 547017 398414 578898
rect 401514 705798 402134 705830
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547017 402134 582618
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 547017 434414 578898
rect 437514 705798 438134 705830
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 460979 632092 461045 632093
rect 460979 632028 460980 632092
rect 461044 632028 461045 632092
rect 460979 632027 461045 632028
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547017 438134 582618
rect 460059 557836 460125 557837
rect 460059 557772 460060 557836
rect 460124 557772 460125 557836
rect 460059 557771 460125 557772
rect 451043 556884 451109 556885
rect 451043 556820 451044 556884
rect 451108 556820 451109 556884
rect 451043 556819 451109 556820
rect 231347 535940 231413 535941
rect 231347 535876 231348 535940
rect 231412 535876 231413 535940
rect 231347 535875 231413 535876
rect 231163 300116 231229 300117
rect 231163 300052 231164 300116
rect 231228 300052 231229 300116
rect 231163 300051 231229 300052
rect 231350 170373 231410 535875
rect 233371 523700 233437 523701
rect 233371 523636 233372 523700
rect 233436 523636 233437 523700
rect 233371 523635 233437 523636
rect 231715 512140 231781 512141
rect 231715 512076 231716 512140
rect 231780 512076 231781 512140
rect 231715 512075 231781 512076
rect 231531 497860 231597 497861
rect 231531 497796 231532 497860
rect 231596 497796 231597 497860
rect 231531 497795 231597 497796
rect 231347 170372 231413 170373
rect 231347 170308 231348 170372
rect 231412 170308 231413 170372
rect 231347 170307 231413 170308
rect 231534 36549 231594 497795
rect 231718 37909 231778 512075
rect 233003 467260 233069 467261
rect 233003 467196 233004 467260
rect 233068 467196 233069 467260
rect 233003 467195 233069 467196
rect 232819 437340 232885 437341
rect 232819 437276 232820 437340
rect 232884 437276 232885 437340
rect 232819 437275 232885 437276
rect 232635 406740 232701 406741
rect 232635 406676 232636 406740
rect 232700 406676 232701 406740
rect 232635 406675 232701 406676
rect 232451 388380 232517 388381
rect 232451 388316 232452 388380
rect 232516 388316 232517 388380
rect 232451 388315 232517 388316
rect 232454 318205 232514 388315
rect 232451 318204 232517 318205
rect 232451 318140 232452 318204
rect 232516 318140 232517 318204
rect 232451 318139 232517 318140
rect 232638 316845 232698 406675
rect 232822 337381 232882 437275
rect 232819 337380 232885 337381
rect 232819 337316 232820 337380
rect 232884 337316 232885 337380
rect 232819 337315 232885 337316
rect 232635 316844 232701 316845
rect 232635 316780 232636 316844
rect 232700 316780 232701 316844
rect 232635 316779 232701 316780
rect 233006 293181 233066 467195
rect 233187 447540 233253 447541
rect 233187 447476 233188 447540
rect 233252 447476 233253 447540
rect 233187 447475 233253 447476
rect 233190 331805 233250 447475
rect 233187 331804 233253 331805
rect 233187 331740 233188 331804
rect 233252 331740 233253 331804
rect 233187 331739 233253 331740
rect 233374 329221 233434 523635
rect 233739 503980 233805 503981
rect 233739 503916 233740 503980
rect 233804 503916 233805 503980
rect 233739 503915 233805 503916
rect 233555 469980 233621 469981
rect 233555 469916 233556 469980
rect 233620 469916 233621 469980
rect 233555 469915 233621 469916
rect 233371 329220 233437 329221
rect 233371 329156 233372 329220
rect 233436 329156 233437 329220
rect 233371 329155 233437 329156
rect 233003 293180 233069 293181
rect 233003 293116 233004 293180
rect 233068 293116 233069 293180
rect 233003 293115 233069 293116
rect 233558 258773 233618 469915
rect 233555 258772 233621 258773
rect 233555 258708 233556 258772
rect 233620 258708 233621 258772
rect 233555 258707 233621 258708
rect 233742 111893 233802 503915
rect 235027 427820 235093 427821
rect 235027 427756 235028 427820
rect 235092 427756 235093 427820
rect 235027 427755 235093 427756
rect 235030 327861 235090 427755
rect 450859 404020 450925 404021
rect 450859 403956 450860 404020
rect 450924 403956 450925 404020
rect 450859 403955 450925 403956
rect 450862 393330 450922 403955
rect 450310 393270 450922 393330
rect 235211 387020 235277 387021
rect 235211 386956 235212 387020
rect 235276 386956 235277 387020
rect 235211 386955 235277 386956
rect 235027 327860 235093 327861
rect 235027 327796 235028 327860
rect 235092 327796 235093 327860
rect 235027 327795 235093 327796
rect 235214 318069 235274 386955
rect 235395 358460 235461 358461
rect 235395 358396 235396 358460
rect 235460 358396 235461 358460
rect 235395 358395 235461 358396
rect 235398 336701 235458 358395
rect 328499 339964 328565 339965
rect 328499 339900 328500 339964
rect 328564 339900 328565 339964
rect 328499 339899 328565 339900
rect 391795 339964 391861 339965
rect 391795 339900 391796 339964
rect 391860 339900 391861 339964
rect 391795 339899 391861 339900
rect 237419 339828 237485 339829
rect 237419 339764 237420 339828
rect 237484 339764 237485 339828
rect 237419 339763 237485 339764
rect 237235 339012 237301 339013
rect 237235 338948 237236 339012
rect 237300 338948 237301 339012
rect 237235 338947 237301 338948
rect 237238 337925 237298 338947
rect 237235 337924 237301 337925
rect 237235 337860 237236 337924
rect 237300 337860 237301 337924
rect 237235 337859 237301 337860
rect 237422 337517 237482 339763
rect 262811 338876 262877 338877
rect 262811 338812 262812 338876
rect 262876 338812 262877 338876
rect 262811 338811 262877 338812
rect 237419 337516 237485 337517
rect 237419 337452 237420 337516
rect 237484 337452 237485 337516
rect 237419 337451 237485 337452
rect 235395 336700 235461 336701
rect 235395 336636 235396 336700
rect 235460 336636 235461 336700
rect 235395 336635 235461 336636
rect 253794 327454 254414 338423
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 235211 318068 235277 318069
rect 235211 318004 235212 318068
rect 235276 318004 235277 318068
rect 235211 318003 235277 318004
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 233739 111892 233805 111893
rect 233739 111828 233740 111892
rect 233804 111828 233805 111892
rect 233739 111827 233805 111828
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 231715 37908 231781 37909
rect 231715 37844 231716 37908
rect 231780 37844 231781 37908
rect 231715 37843 231781 37844
rect 231531 36548 231597 36549
rect 231531 36484 231532 36548
rect 231596 36484 231597 36548
rect 231531 36483 231597 36484
rect 229691 3908 229757 3909
rect 229691 3844 229692 3908
rect 229756 3844 229757 3908
rect 229691 3843 229757 3844
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -1894 222134 -1862
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 331174 258134 338423
rect 262814 338197 262874 338811
rect 269251 338740 269317 338741
rect 269251 338676 269252 338740
rect 269316 338676 269317 338740
rect 269251 338675 269317 338676
rect 269254 338197 269314 338675
rect 262811 338196 262877 338197
rect 262811 338132 262812 338196
rect 262876 338132 262877 338196
rect 262811 338131 262877 338132
rect 269251 338196 269317 338197
rect 269251 338132 269252 338196
rect 269316 338132 269317 338196
rect 269251 338131 269317 338132
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -1894 258134 -1862
rect 289794 327454 290414 338423
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 331174 294134 338423
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -1894 294134 -1862
rect 325794 327454 326414 338423
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 328502 3229 328562 339899
rect 379651 338740 379717 338741
rect 379651 338676 379652 338740
rect 379716 338676 379717 338740
rect 379651 338675 379717 338676
rect 329514 331174 330134 338423
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 325794 3134 326414 3218
rect 328499 3228 328565 3229
rect 328499 3164 328500 3228
rect 328564 3164 328565 3228
rect 328499 3163 328565 3164
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -1894 330134 -1862
rect 361794 327454 362414 338423
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 331174 366134 338423
rect 379654 338197 379714 338675
rect 379651 338196 379717 338197
rect 379651 338132 379652 338196
rect 379716 338132 379717 338196
rect 379651 338131 379717 338132
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 391798 3501 391858 339899
rect 450123 339828 450189 339829
rect 450123 339764 450124 339828
rect 450188 339764 450189 339828
rect 450123 339763 450189 339764
rect 447731 339692 447797 339693
rect 447731 339628 447732 339692
rect 447796 339628 447797 339692
rect 447731 339627 447797 339628
rect 412403 339012 412469 339013
rect 412403 338948 412404 339012
rect 412468 338948 412469 339012
rect 412403 338947 412469 338948
rect 398971 338876 399037 338877
rect 398971 338812 398972 338876
rect 399036 338812 399037 338876
rect 398971 338811 399037 338812
rect 397794 327454 398414 338423
rect 398974 338197 399034 338811
rect 398971 338196 399037 338197
rect 398971 338132 398972 338196
rect 399036 338132 399037 338196
rect 398971 338131 399037 338132
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 391795 3500 391861 3501
rect 391795 3436 391796 3500
rect 391860 3436 391861 3500
rect 391795 3435 391861 3436
rect 397794 3454 398414 38898
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -1894 366134 -1862
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 331174 402134 338423
rect 412406 338197 412466 338947
rect 412403 338196 412469 338197
rect 412403 338132 412404 338196
rect 412468 338132 412469 338196
rect 412403 338131 412469 338132
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -1894 402134 -1862
rect 433794 327454 434414 338423
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 331174 438134 338423
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 447734 4045 447794 339627
rect 450126 334117 450186 339763
rect 450123 334116 450189 334117
rect 450123 334052 450124 334116
rect 450188 334052 450189 334116
rect 450123 334051 450189 334052
rect 450310 320789 450370 393270
rect 450859 341460 450925 341461
rect 450859 341396 450860 341460
rect 450924 341396 450925 341460
rect 450859 341395 450925 341396
rect 450862 335370 450922 341395
rect 451046 339965 451106 556819
rect 458403 552940 458469 552941
rect 458403 552876 458404 552940
rect 458468 552876 458469 552940
rect 458403 552875 458469 552876
rect 455643 551580 455709 551581
rect 455643 551516 455644 551580
rect 455708 551516 455709 551580
rect 455643 551515 455709 551516
rect 452883 539340 452949 539341
rect 452883 539276 452884 539340
rect 452948 539276 452949 539340
rect 452883 539275 452949 539276
rect 451411 493780 451477 493781
rect 451411 493716 451412 493780
rect 451476 493716 451477 493780
rect 451411 493715 451477 493716
rect 451043 339964 451109 339965
rect 451043 339900 451044 339964
rect 451108 339900 451109 339964
rect 451043 339899 451109 339900
rect 450494 335310 450922 335370
rect 450307 320788 450373 320789
rect 450307 320724 450308 320788
rect 450372 320724 450373 320788
rect 450307 320723 450373 320724
rect 450494 6493 450554 335310
rect 451414 323645 451474 493715
rect 452699 410820 452765 410821
rect 452699 410756 452700 410820
rect 452764 410756 452765 410820
rect 452699 410755 452765 410756
rect 451963 410004 452029 410005
rect 451963 409940 451964 410004
rect 452028 409940 452029 410004
rect 451963 409939 452029 409940
rect 451411 323644 451477 323645
rect 451411 323580 451412 323644
rect 451476 323580 451477 323644
rect 451411 323579 451477 323580
rect 450491 6492 450557 6493
rect 450491 6428 450492 6492
rect 450556 6428 450557 6492
rect 450491 6427 450557 6428
rect 447731 4044 447797 4045
rect 447731 3980 447732 4044
rect 447796 3980 447797 4044
rect 447731 3979 447797 3980
rect 451966 3909 452026 409939
rect 452702 15877 452762 410755
rect 452886 314125 452946 539275
rect 454171 497180 454237 497181
rect 454171 497116 454172 497180
rect 454236 497116 454237 497180
rect 454171 497115 454237 497116
rect 454174 451290 454234 497115
rect 455459 461820 455525 461821
rect 455459 461756 455460 461820
rect 455524 461756 455525 461820
rect 455459 461755 455525 461756
rect 453990 451230 454234 451290
rect 453067 398580 453133 398581
rect 453067 398516 453068 398580
rect 453132 398516 453133 398580
rect 453067 398515 453133 398516
rect 452883 314124 452949 314125
rect 452883 314060 452884 314124
rect 452948 314060 452949 314124
rect 452883 314059 452949 314060
rect 453070 308413 453130 398515
rect 453251 351660 453317 351661
rect 453251 351596 453252 351660
rect 453316 351596 453317 351660
rect 453251 351595 453317 351596
rect 453254 312493 453314 351595
rect 453251 312492 453317 312493
rect 453251 312428 453252 312492
rect 453316 312428 453317 312492
rect 453251 312427 453317 312428
rect 453067 308412 453133 308413
rect 453067 308348 453068 308412
rect 453132 308348 453133 308412
rect 453067 308347 453133 308348
rect 453990 161490 454050 451230
rect 454355 448900 454421 448901
rect 454355 448836 454356 448900
rect 454420 448836 454421 448900
rect 454355 448835 454421 448836
rect 454171 446180 454237 446181
rect 454171 446116 454172 446180
rect 454236 446116 454237 446180
rect 454171 446115 454237 446116
rect 454174 166293 454234 446115
rect 454358 301477 454418 448835
rect 454539 422380 454605 422381
rect 454539 422316 454540 422380
rect 454604 422316 454605 422380
rect 454539 422315 454605 422316
rect 454542 311133 454602 422315
rect 454539 311132 454605 311133
rect 454539 311068 454540 311132
rect 454604 311068 454605 311132
rect 454539 311067 454605 311068
rect 454355 301476 454421 301477
rect 454355 301412 454356 301476
rect 454420 301412 454421 301476
rect 454355 301411 454421 301412
rect 454171 166292 454237 166293
rect 454171 166228 454172 166292
rect 454236 166228 454237 166292
rect 454171 166227 454237 166228
rect 453990 161430 454234 161490
rect 452699 15876 452765 15877
rect 452699 15812 452700 15876
rect 452764 15812 452765 15876
rect 452699 15811 452765 15812
rect 454174 11661 454234 161430
rect 455462 112437 455522 461755
rect 455646 323781 455706 551515
rect 458219 529140 458285 529141
rect 458219 529076 458220 529140
rect 458284 529076 458285 529140
rect 458219 529075 458285 529076
rect 456747 523700 456813 523701
rect 456747 523636 456748 523700
rect 456812 523636 456813 523700
rect 456747 523635 456813 523636
rect 456011 415580 456077 415581
rect 456011 415516 456012 415580
rect 456076 415516 456077 415580
rect 456011 415515 456077 415516
rect 455827 412180 455893 412181
rect 455827 412116 455828 412180
rect 455892 412116 455893 412180
rect 455827 412115 455893 412116
rect 455643 323780 455709 323781
rect 455643 323716 455644 323780
rect 455708 323716 455709 323780
rect 455643 323715 455709 323716
rect 455830 296037 455890 412115
rect 456014 316709 456074 415515
rect 456011 316708 456077 316709
rect 456011 316644 456012 316708
rect 456076 316644 456077 316708
rect 456011 316643 456077 316644
rect 455827 296036 455893 296037
rect 455827 295972 455828 296036
rect 455892 295972 455893 296036
rect 455827 295971 455893 295972
rect 456750 251837 456810 523635
rect 456931 505340 456997 505341
rect 456931 505276 456932 505340
rect 456996 505276 456997 505340
rect 456931 505275 456997 505276
rect 456934 315349 456994 505275
rect 457115 443460 457181 443461
rect 457115 443396 457116 443460
rect 457180 443396 457181 443460
rect 457115 443395 457181 443396
rect 457118 327725 457178 443395
rect 457299 433260 457365 433261
rect 457299 433196 457300 433260
rect 457364 433196 457365 433260
rect 457299 433195 457365 433196
rect 457115 327724 457181 327725
rect 457115 327660 457116 327724
rect 457180 327660 457181 327724
rect 457115 327659 457181 327660
rect 457302 320925 457362 433195
rect 457299 320924 457365 320925
rect 457299 320860 457300 320924
rect 457364 320860 457365 320924
rect 457299 320859 457365 320860
rect 456931 315348 456997 315349
rect 456931 315284 456932 315348
rect 456996 315284 456997 315348
rect 456931 315283 456997 315284
rect 458222 283525 458282 529075
rect 458406 309773 458466 552875
rect 458587 548860 458653 548861
rect 458587 548796 458588 548860
rect 458652 548796 458653 548860
rect 458587 548795 458653 548796
rect 458590 313989 458650 548795
rect 458771 501260 458837 501261
rect 458771 501196 458772 501260
rect 458836 501196 458837 501260
rect 458771 501195 458837 501196
rect 458774 322149 458834 501195
rect 459507 484260 459573 484261
rect 459507 484196 459508 484260
rect 459572 484196 459573 484260
rect 459507 484195 459573 484196
rect 459510 336157 459570 484195
rect 459507 336156 459573 336157
rect 459507 336092 459508 336156
rect 459572 336092 459573 336156
rect 459507 336091 459573 336092
rect 458771 322148 458837 322149
rect 458771 322084 458772 322148
rect 458836 322084 458837 322148
rect 458771 322083 458837 322084
rect 458587 313988 458653 313989
rect 458587 313924 458588 313988
rect 458652 313924 458653 313988
rect 458587 313923 458653 313924
rect 458403 309772 458469 309773
rect 458403 309708 458404 309772
rect 458468 309708 458469 309772
rect 458403 309707 458469 309708
rect 458219 283524 458285 283525
rect 458219 283460 458220 283524
rect 458284 283460 458285 283524
rect 458219 283459 458285 283460
rect 456747 251836 456813 251837
rect 456747 251772 456748 251836
rect 456812 251772 456813 251836
rect 456747 251771 456813 251772
rect 455459 112436 455525 112437
rect 455459 112372 455460 112436
rect 455524 112372 455525 112436
rect 455459 112371 455525 112372
rect 454171 11660 454237 11661
rect 454171 11596 454172 11660
rect 454236 11596 454237 11660
rect 454171 11595 454237 11596
rect 451963 3908 452029 3909
rect 451963 3844 451964 3908
rect 452028 3844 452029 3908
rect 451963 3843 452029 3844
rect 460062 3501 460122 557771
rect 460243 556612 460309 556613
rect 460243 556548 460244 556612
rect 460308 556548 460309 556612
rect 460243 556547 460309 556548
rect 460059 3500 460125 3501
rect 460059 3436 460060 3500
rect 460124 3436 460125 3500
rect 460059 3435 460125 3436
rect 460246 3365 460306 556547
rect 460982 360229 461042 632027
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 461163 559060 461229 559061
rect 461163 558996 461164 559060
rect 461228 558996 461229 559060
rect 461163 558995 461229 558996
rect 460979 360228 461045 360229
rect 460979 360164 460980 360228
rect 461044 360164 461045 360228
rect 460979 360163 461045 360164
rect 461166 336565 461226 558995
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 463739 510644 463805 510645
rect 463739 510580 463740 510644
rect 463804 510580 463805 510644
rect 463739 510579 463805 510580
rect 461347 506564 461413 506565
rect 461347 506500 461348 506564
rect 461412 506500 461413 506564
rect 461347 506499 461413 506500
rect 461163 336564 461229 336565
rect 461163 336500 461164 336564
rect 461228 336500 461229 336564
rect 461163 336499 461229 336500
rect 461350 336293 461410 506499
rect 462267 441692 462333 441693
rect 462267 441628 462268 441692
rect 462332 441628 462333 441692
rect 462267 441627 462333 441628
rect 461347 336292 461413 336293
rect 461347 336228 461348 336292
rect 461412 336228 461413 336292
rect 461347 336227 461413 336228
rect 462270 334661 462330 441627
rect 462267 334660 462333 334661
rect 462267 334596 462268 334660
rect 462332 334596 462333 334660
rect 462267 334595 462333 334596
rect 463742 333573 463802 510579
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 463739 333572 463805 333573
rect 463739 333508 463740 333572
rect 463804 333508 463805 333572
rect 463739 333507 463805 333508
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 460243 3364 460309 3365
rect 460243 3300 460244 3364
rect 460308 3300 460309 3364
rect 460243 3299 460309 3300
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -1894 438134 -1862
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 705798 474134 705830
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -1894 474134 -1862
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 705798 510134 705830
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -1894 510134 -1862
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 705798 546134 705830
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -1894 546134 -1862
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 705798 582134 705830
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -1894 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
<< via4 >>
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
<< metal5 >>
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -2966 691174 586890 691206
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect -2966 690854 586890 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect -2966 690586 586890 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -2966 655174 586890 655206
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect -2966 654854 586890 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect -2966 654586 586890 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -2966 619174 586890 619206
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect -2966 618854 586890 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect -2966 618586 586890 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -2966 583174 586890 583206
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect -2966 582854 586890 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect -2966 582586 586890 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -2966 547174 586890 547206
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect -2966 546854 586890 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect -2966 546586 586890 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -2966 511174 234820 511206
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 234820 511174
rect -2966 510854 234820 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 234820 510854
rect -2966 510586 234820 510618
rect 375572 511174 586890 511206
rect 375572 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 375572 510854 586890 510938
rect 375572 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 375572 510586 586890 510618
rect -2966 507454 234820 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 234820 507454
rect -2966 507134 234820 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 234820 507134
rect -2966 506866 234820 506898
rect 375572 507454 586890 507486
rect 375572 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect 375572 507134 586890 507218
rect 375572 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect 375572 506866 586890 506898
rect -2966 475174 234820 475206
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 234820 475174
rect -2966 474854 234820 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 234820 474854
rect -2966 474586 234820 474618
rect 375572 475174 586890 475206
rect 375572 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 375572 474854 586890 474938
rect 375572 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 375572 474586 586890 474618
rect -2966 471454 234820 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 234820 471454
rect -2966 471134 234820 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 234820 471134
rect -2966 470866 234820 470898
rect 375572 471454 586890 471486
rect 375572 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect 375572 471134 586890 471218
rect 375572 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect 375572 470866 586890 470898
rect -2966 439174 234820 439206
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 234820 439174
rect -2966 438854 234820 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 234820 438854
rect -2966 438586 234820 438618
rect 375572 439174 586890 439206
rect 375572 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 375572 438854 586890 438938
rect 375572 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 375572 438586 586890 438618
rect -2966 435454 234820 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 234820 435454
rect -2966 435134 234820 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 234820 435134
rect -2966 434866 234820 434898
rect 375572 435454 586890 435486
rect 375572 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect 375572 435134 586890 435218
rect 375572 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect 375572 434866 586890 434898
rect -2966 403174 234820 403206
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 234820 403174
rect -2966 402854 234820 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 234820 402854
rect -2966 402586 234820 402618
rect 375572 403174 586890 403206
rect 375572 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 375572 402854 586890 402938
rect 375572 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 375572 402586 586890 402618
rect -2966 399454 234820 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 234820 399454
rect -2966 399134 234820 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 234820 399134
rect -2966 398866 234820 398898
rect 375572 399454 586890 399486
rect 375572 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect 375572 399134 586890 399218
rect 375572 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect 375572 398866 586890 398898
rect -2966 367174 234820 367206
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 234820 367174
rect -2966 366854 234820 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 234820 366854
rect -2966 366586 234820 366618
rect 375572 367174 586890 367206
rect 375572 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 375572 366854 586890 366938
rect 375572 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 375572 366586 586890 366618
rect -2966 363454 234820 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 234820 363454
rect -2966 363134 234820 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 234820 363134
rect -2966 362866 234820 362898
rect 375572 363454 586890 363486
rect 375572 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect 375572 363134 586890 363218
rect 375572 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect 375572 362866 586890 362898
rect -2966 331174 586890 331206
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect -2966 330854 586890 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect -2966 330586 586890 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -2966 295174 586890 295206
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect -2966 294854 586890 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect -2966 294586 586890 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -2966 259174 586890 259206
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect -2966 258854 586890 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect -2966 258586 586890 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -2966 223174 586890 223206
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect -2966 222854 586890 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect -2966 222586 586890 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -2966 187174 586890 187206
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect -2966 186854 586890 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect -2966 186586 586890 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -2966 151174 586890 151206
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect -2966 150854 586890 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect -2966 150586 586890 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -2966 115174 586890 115206
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect -2966 114854 586890 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect -2966 114586 586890 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -2966 79174 586890 79206
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect -2966 78854 586890 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect -2966 78586 586890 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -2966 43174 586890 43206
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect -2966 42854 586890 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect -2966 42586 586890 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -2966 7174 586890 7206
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect -2966 6854 586890 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect -2966 6586 586890 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
use soc_now_caravel_top  mprj
timestamp 0
transform 1 0 235000 0 1 338000
box -1076 -4 217552 218628
<< labels >>
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5514 -1894 6134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 41514 -1894 42134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 77514 -1894 78134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 113514 -1894 114134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 149514 -1894 150134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 185514 -1894 186134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 221514 -1894 222134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 257514 -1894 258134 338423 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 257514 547017 258134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 293514 -1894 294134 338423 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 293514 547017 294134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 329514 -1894 330134 338423 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 329514 547017 330134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 365514 -1894 366134 338423 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 365514 547017 366134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 401514 -1894 402134 338423 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 401514 547017 402134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 437514 -1894 438134 338423 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 437514 547017 438134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 473514 -1894 474134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 509514 -1894 510134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 545514 -1894 546134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 581514 -1894 582134 705830 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 6586 586890 7206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 42586 586890 43206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 78586 586890 79206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 114586 586890 115206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 150586 586890 151206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 186586 586890 187206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 222586 586890 223206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 258586 586890 259206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 294586 586890 295206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 330586 586890 331206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 366586 234820 367206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 402586 234820 403206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 438586 234820 439206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 474586 234820 475206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 510586 234820 511206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 546586 586890 547206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 582586 586890 583206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 618586 586890 619206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 654586 586890 655206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 690586 586890 691206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 375572 366586 586890 367206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 375572 402586 586890 403206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 375572 438586 586890 439206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 375572 474586 586890 475206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 375572 510586 586890 511206 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 1794 -1894 2414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 37794 -1894 38414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 73794 -1894 74414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 109794 -1894 110414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 145794 -1894 146414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 181794 -1894 182414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 217794 -1894 218414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 253794 -1894 254414 338423 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 253794 547017 254414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 289794 -1894 290414 338423 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 289794 547017 290414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 325794 -1894 326414 338423 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 325794 547017 326414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 361794 -1894 362414 338423 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 361794 547017 362414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 397794 -1894 398414 338423 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 397794 547017 398414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 433794 -1894 434414 338423 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 433794 547017 434414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 469794 -1894 470414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 505794 -1894 506414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 541794 -1894 542414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 577794 -1894 578414 705830 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 2866 586890 3486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 38866 586890 39486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 74866 586890 75486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 110866 586890 111486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 146866 586890 147486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 182866 586890 183486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 218866 586890 219486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 254866 586890 255486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 290866 586890 291486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 326866 586890 327486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 362866 234820 363486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 398866 234820 399486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 434866 234820 435486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 470866 234820 471486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 506866 234820 507486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 542866 586890 543486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 578866 586890 579486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 614866 586890 615486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 650866 586890 651486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 686866 586890 687486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 375572 362866 586890 363486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 375572 398866 586890 399486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 375572 434866 586890 435486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 375572 470866 586890 471486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 375572 506866 586890 507486 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 2 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 3 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 4 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 5 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 6 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 7 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 8 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 9 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 10 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 11 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 12 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 13 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 14 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 15 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 16 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 17 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 18 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 19 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 20 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 21 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 22 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 23 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 24 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 25 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 26 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 27 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 28 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 29 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 30 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 31 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 32 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 33 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 34 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 35 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 36 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 37 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 38 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 39 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 40 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 41 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 42 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 43 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 44 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 45 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 46 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 47 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 48 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 49 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 50 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 51 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 52 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 53 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 54 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 55 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 56 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 57 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 58 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 59 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 60 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 61 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 62 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 63 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 64 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 65 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 66 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 67 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 68 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 69 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 70 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 71 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 72 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 73 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 74 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 75 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 76 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 77 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 78 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 79 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 80 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 81 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 82 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 83 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 84 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 85 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 86 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 87 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 88 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 89 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 90 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 91 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 92 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 93 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 94 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 95 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 96 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 97 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 98 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 99 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 100 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 101 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 102 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 103 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 104 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 105 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 106 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 107 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 108 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 109 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 110 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 111 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 112 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 113 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 114 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 115 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 116 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 117 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 118 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 119 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 120 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 121 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 122 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 123 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 124 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 125 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 126 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 127 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 128 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 129 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 130 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 131 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 132 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 133 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 134 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 135 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 136 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 137 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 138 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 139 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 140 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 141 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 142 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 143 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 144 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 145 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 146 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 147 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 148 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 149 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 150 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 151 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 152 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 153 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 154 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 155 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 156 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 157 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 158 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 159 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 160 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 161 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 162 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 163 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 164 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 165 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 166 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 167 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 168 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 169 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 170 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 171 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 172 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 173 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 174 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 175 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 176 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 177 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 178 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 179 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 180 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 181 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 182 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 183 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 184 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 185 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 186 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 187 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 188 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 189 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 190 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 191 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 192 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 193 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 194 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 195 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 196 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 197 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 198 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 199 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 200 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 201 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 202 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 203 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 204 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 205 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 206 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 207 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 208 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 209 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 210 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 211 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 212 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 213 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 214 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 215 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 216 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 217 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 218 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 219 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 220 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 221 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 222 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 223 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 224 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 225 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 226 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 227 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 228 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 229 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 230 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 231 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 232 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 233 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 234 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 235 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 236 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 237 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 238 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 239 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 240 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 241 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 242 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 243 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 244 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 245 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 246 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 247 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 248 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 249 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 250 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 251 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 252 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 253 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 254 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 255 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 256 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 257 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 258 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 259 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 260 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 261 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 262 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 263 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 264 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 265 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 266 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 267 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 268 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 269 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 270 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 271 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 272 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 273 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 274 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 275 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 276 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 277 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 278 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 279 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 280 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 281 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 282 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 283 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 284 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 285 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 286 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 287 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 288 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 289 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 290 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 291 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 292 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 293 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 294 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 295 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 296 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 297 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 298 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 299 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 300 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 301 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 302 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 303 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 304 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 305 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 306 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 307 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 308 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 309 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 310 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 311 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 312 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 313 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 314 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 315 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 316 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 317 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 318 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 319 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 320 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 321 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 322 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 323 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 324 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 325 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 326 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 327 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 328 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 329 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 330 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 331 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 332 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 333 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 334 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 335 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 336 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 337 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 338 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 339 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 340 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 341 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 342 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 343 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 344 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 345 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 346 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 347 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 348 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 349 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 350 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 351 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 352 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 353 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 354 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 355 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 356 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 357 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 358 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 359 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 360 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 361 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 362 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 363 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 364 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 365 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 366 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 367 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 368 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 369 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 370 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 371 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 372 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 373 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 374 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 375 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 376 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 377 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 378 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 379 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 380 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 381 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 382 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 383 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 384 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 385 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 386 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 387 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 388 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 389 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 390 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 391 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 392 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 393 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 394 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 395 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 396 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 397 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 398 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 399 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 400 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 401 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 402 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 403 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 404 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 405 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 406 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 407 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 408 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 409 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 410 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 411 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 412 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 413 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 414 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 415 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 416 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 417 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 418 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 419 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 420 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 421 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 422 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 423 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 424 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 425 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 426 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 427 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 428 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 429 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 430 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 431 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 432 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 433 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 434 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 435 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 436 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 437 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 438 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 439 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 440 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 441 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 442 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 443 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 444 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 445 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 446 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 447 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 448 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 449 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 450 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 451 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 452 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 453 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 454 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 455 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 456 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 457 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 458 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 459 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 460 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 461 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 462 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 463 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 464 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 465 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 466 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 467 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 468 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 469 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 470 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 471 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 472 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 473 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 474 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 475 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 476 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 477 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 478 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 479 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 480 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 481 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 482 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 483 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 484 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 485 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 486 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 487 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 488 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 489 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 490 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 491 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 492 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 493 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 494 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 495 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 496 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 497 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 498 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 499 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 500 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 501 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 502 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 503 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 504 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 505 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 506 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 507 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 508 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 509 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 510 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 511 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 512 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 513 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 514 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 515 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 516 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 517 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 518 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 519 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 520 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 521 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 522 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 523 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 524 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 525 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 526 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 527 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 528 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 529 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 530 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 531 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 532 nsew signal tristate
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 533 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 534 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 535 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 536 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 537 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 538 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 539 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 540 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 541 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 542 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 543 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 544 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 545 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 546 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 547 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 548 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 549 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 550 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 551 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 552 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 553 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 554 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 555 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 556 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 557 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 558 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 559 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 560 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 561 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 562 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 563 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 564 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 565 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 566 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 567 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 568 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 569 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 570 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 571 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 572 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 573 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 574 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 575 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 576 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 577 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 578 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 579 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 580 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 581 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 582 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 583 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 584 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 585 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 586 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 587 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 588 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 589 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 590 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 591 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 592 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 593 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 594 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 595 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 596 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 597 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 598 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 599 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 600 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 601 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 602 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 603 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 604 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 605 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 606 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 607 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 608 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 609 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 610 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 611 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 612 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 613 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 614 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 615 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 616 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 617 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 618 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 619 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 620 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 621 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 622 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 623 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 624 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 625 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 626 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 627 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 628 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 629 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 630 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 631 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 632 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 633 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 634 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 635 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 636 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 637 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 638 nsew signal input
rlabel metal5 481231 510896 481231 510896 0 VGND
rlabel metal5 481231 507176 481231 507176 0 VPWR
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal2 232070 351101 232070 351101 0 io_in[10]
rlabel metal2 541650 467840 541650 467840 0 io_in[11]
rlabel metal2 579830 563703 579830 563703 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel metal2 580198 670735 580198 670735 0 io_in[14]
rlabel metal2 252234 556580 252234 556580 0 io_in[15]
rlabel metal3 234792 547468 234792 547468 0 io_in[16]
rlabel metal2 429456 703596 429456 703596 0 io_in[17]
rlabel metal3 234102 495108 234102 495108 0 io_in[18]
rlabel metal2 306974 556580 306974 556580 0 io_in[19]
rlabel metal2 507150 303654 507150 303654 0 io_in[1]
rlabel metal2 234830 703596 234830 703596 0 io_in[20]
rlabel metal3 452356 508028 452356 508028 0 io_in[21]
rlabel metal3 452724 385628 452724 385628 0 io_in[22]
rlabel metal2 40204 703596 40204 703596 0 io_in[23]
rlabel metal3 1878 684284 1878 684284 0 io_in[24]
rlabel metal4 461012 496128 461012 496128 0 io_in[25]
rlabel metal3 1832 579972 1832 579972 0 io_in[26]
rlabel metal3 1832 527884 1832 527884 0 io_in[27]
rlabel metal3 1832 475660 1832 475660 0 io_in[28]
rlabel metal3 1740 423572 1740 423572 0 io_in[29]
rlabel metal2 232070 526099 232070 526099 0 io_in[2]
rlabel metal3 1924 371348 1924 371348 0 io_in[30]
rlabel metal3 1924 319260 1924 319260 0 io_in[31]
rlabel metal3 1924 267172 1924 267172 0 io_in[32]
rlabel metal3 1832 214948 1832 214948 0 io_in[33]
rlabel metal3 1786 162860 1786 162860 0 io_in[34]
rlabel metal3 1878 110636 1878 110636 0 io_in[35]
rlabel metal3 1878 71604 1878 71604 0 io_in[36]
rlabel metal3 1924 32436 1924 32436 0 io_in[37]
rlabel metal2 423276 556580 423276 556580 0 io_in[3]
rlabel metal2 232070 537047 232070 537047 0 io_in[4]
rlabel metal2 580014 206329 580014 206329 0 io_in[5]
rlabel metal2 232070 441847 232070 441847 0 io_in[6]
rlabel metal2 468602 426428 468602 426428 0 io_in[7]
rlabel metal3 582092 351900 582092 351900 0 io_in[8]
rlabel metal2 580198 404651 580198 404651 0 io_in[9]
rlabel via2 580198 33099 580198 33099 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal2 275156 338028 275156 338028 0 io_oeb[11]
rlabel metal1 450570 336736 450570 336736 0 io_oeb[12]
rlabel metal2 580198 643569 580198 643569 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal2 232990 504356 232990 504356 0 io_oeb[15]
rlabel metal1 462024 699686 462024 699686 0 io_oeb[16]
rlabel metal3 452724 347548 452724 347548 0 io_oeb[17]
rlabel metal2 256098 556580 256098 556580 0 io_oeb[18]
rlabel metal1 351900 700366 351900 700366 0 io_oeb[19]
rlabel metal2 232070 539801 232070 539801 0 io_oeb[1]
rlabel metal2 231978 344913 231978 344913 0 io_oeb[20]
rlabel metal2 137862 702008 137862 702008 0 io_oeb[21]
rlabel metal1 72404 703018 72404 703018 0 io_oeb[22]
rlabel metal1 69966 700366 69966 700366 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal3 1878 606084 1878 606084 0 io_oeb[25]
rlabel metal2 232070 408255 232070 408255 0 io_oeb[26]
rlabel metal3 1786 501772 1786 501772 0 io_oeb[27]
rlabel metal3 1832 449548 1832 449548 0 io_oeb[28]
rlabel metal3 1832 397460 1832 397460 0 io_oeb[29]
rlabel metal3 234401 503948 234401 503948 0 io_oeb[2]
rlabel metal3 1832 345372 1832 345372 0 io_oeb[30]
rlabel metal3 1924 293148 1924 293148 0 io_oeb[31]
rlabel metal3 1878 241060 1878 241060 0 io_oeb[32]
rlabel metal3 1878 188836 1878 188836 0 io_oeb[33]
rlabel metal2 348190 556580 348190 556580 0 io_oeb[34]
rlabel metal3 1740 84660 1740 84660 0 io_oeb[35]
rlabel metal3 1878 45492 1878 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580014 152915 580014 152915 0 io_oeb[3]
rlabel metal2 580198 192831 580198 192831 0 io_oeb[4]
rlabel metal3 581954 232356 581954 232356 0 io_oeb[5]
rlabel metal2 580198 272697 580198 272697 0 io_oeb[6]
rlabel metal2 330112 338028 330112 338028 0 io_oeb[7]
rlabel metal2 253260 338028 253260 338028 0 io_oeb[8]
rlabel metal2 580198 430729 580198 430729 0 io_oeb[9]
rlabel metal2 580014 20213 580014 20213 0 io_out[0]
rlabel metal2 424994 337059 424994 337059 0 io_out[10]
rlabel metal2 232070 368577 232070 368577 0 io_out[11]
rlabel metal3 234608 484228 234608 484228 0 io_out[12]
rlabel metal2 237514 556580 237514 556580 0 io_out[13]
rlabel metal2 580198 683519 580198 683519 0 io_out[14]
rlabel metal2 408082 556580 408082 556580 0 io_out[15]
rlabel metal2 255146 338028 255146 338028 0 io_out[16]
rlabel metal3 234654 468588 234654 468588 0 io_out[17]
rlabel metal3 234700 409428 234700 409428 0 io_out[18]
rlabel metal2 282946 636555 282946 636555 0 io_out[19]
rlabel metal3 234309 469948 234309 469948 0 io_out[1]
rlabel metal2 218546 703596 218546 703596 0 io_out[20]
rlabel metal2 154146 701974 154146 701974 0 io_out[21]
rlabel metal1 158148 700298 158148 700298 0 io_out[22]
rlabel metal2 23828 703596 23828 703596 0 io_out[23]
rlabel metal3 1924 671228 1924 671228 0 io_out[24]
rlabel metal3 1740 619140 1740 619140 0 io_out[25]
rlabel metal3 1878 566916 1878 566916 0 io_out[26]
rlabel metal3 1832 514828 1832 514828 0 io_out[27]
rlabel metal3 1970 462604 1970 462604 0 io_out[28]
rlabel metal3 1832 410516 1832 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal3 1924 358428 1924 358428 0 io_out[30]
rlabel metal3 1924 306204 1924 306204 0 io_out[31]
rlabel metal3 1740 254116 1740 254116 0 io_out[32]
rlabel metal3 1878 201892 1878 201892 0 io_out[33]
rlabel metal3 1878 149804 1878 149804 0 io_out[34]
rlabel metal3 1878 97580 1878 97580 0 io_out[35]
rlabel metal3 475 58548 475 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel via2 580198 139349 580198 139349 0 io_out[3]
rlabel metal2 580198 179265 580198 179265 0 io_out[4]
rlabel metal3 581908 219028 581908 219028 0 io_out[5]
rlabel metal3 234700 405348 234700 405348 0 io_out[6]
rlabel metal2 580198 312647 580198 312647 0 io_out[7]
rlabel metal2 580198 364735 580198 364735 0 io_out[8]
rlabel metal2 579738 418217 579738 418217 0 io_out[9]
rlabel metal2 232070 480879 232070 480879 0 la_data_in[0]
rlabel metal2 480424 16560 480424 16560 0 la_data_in[100]
rlabel metal2 329514 556580 329514 556580 0 la_data_in[101]
rlabel metal2 487409 340 487409 340 0 la_data_in[102]
rlabel metal2 468510 275672 468510 275672 0 la_data_in[103]
rlabel metal3 452724 426428 452724 426428 0 la_data_in[104]
rlabel metal3 234608 401268 234608 401268 0 la_data_in[105]
rlabel metal2 501577 340 501577 340 0 la_data_in[106]
rlabel metal3 234125 447508 234125 447508 0 la_data_in[107]
rlabel metal3 234217 523668 234217 523668 0 la_data_in[108]
rlabel via1 296470 556325 296470 556325 0 la_data_in[109]
rlabel metal2 161322 1894 161322 1894 0 la_data_in[10]
rlabel metal2 331246 163161 331246 163161 0 la_data_in[110]
rlabel metal2 519248 16560 519248 16560 0 la_data_in[111]
rlabel metal2 232070 348347 232070 348347 0 la_data_in[112]
rlabel metal1 271032 330446 271032 330446 0 la_data_in[113]
rlabel metal2 232070 489107 232070 489107 0 la_data_in[114]
rlabel metal2 371266 165949 371266 165949 0 la_data_in[115]
rlabel metal3 452724 546108 452724 546108 0 la_data_in[116]
rlabel metal2 526470 219776 526470 219776 0 la_data_in[117]
rlabel metal2 544410 6722 544410 6722 0 la_data_in[118]
rlabel metal2 543030 243576 543030 243576 0 la_data_in[119]
rlabel metal2 232070 460003 232070 460003 0 la_data_in[11]
rlabel metal2 551257 340 551257 340 0 la_data_in[120]
rlabel metal3 452724 499868 452724 499868 0 la_data_in[121]
rlabel metal2 558072 16560 558072 16560 0 la_data_in[122]
rlabel metal2 562074 3968 562074 3968 0 la_data_in[123]
rlabel metal2 565662 1996 565662 1996 0 la_data_in[124]
rlabel metal2 387474 338028 387474 338028 0 la_data_in[125]
rlabel metal2 572746 1826 572746 1826 0 la_data_in[126]
rlabel metal2 562350 181152 562350 181152 0 la_data_in[127]
rlabel via2 232070 425085 232070 425085 0 la_data_in[12]
rlabel metal2 171580 16560 171580 16560 0 la_data_in[13]
rlabel metal2 175398 16560 175398 16560 0 la_data_in[14]
rlabel metal2 179078 2183 179078 2183 0 la_data_in[15]
rlabel metal4 461380 421396 461380 421396 0 la_data_in[16]
rlabel metal3 450409 337620 450409 337620 0 la_data_in[17]
rlabel metal2 448546 315651 448546 315651 0 la_data_in[18]
rlabel metal2 193246 1911 193246 1911 0 la_data_in[19]
rlabel metal2 232070 524739 232070 524739 0 la_data_in[1]
rlabel metal2 232070 383979 232070 383979 0 la_data_in[20]
rlabel metal2 462346 347446 462346 347446 0 la_data_in[21]
rlabel metal2 232070 470951 232070 470951 0 la_data_in[22]
rlabel metal2 248584 556672 248584 556672 0 la_data_in[23]
rlabel metal2 211002 4988 211002 4988 0 la_data_in[24]
rlabel metal2 214222 16560 214222 16560 0 la_data_in[25]
rlabel metal2 218086 278518 218086 278518 0 la_data_in[26]
rlabel metal2 327106 163161 327106 163161 0 la_data_in[27]
rlabel metal3 452724 444788 452724 444788 0 la_data_in[28]
rlabel metal2 228521 340 228521 340 0 la_data_in[29]
rlabel metal2 132756 16560 132756 16560 0 la_data_in[2]
rlabel metal2 232063 340 232063 340 0 la_data_in[30]
rlabel metal2 235842 6722 235842 6722 0 la_data_in[31]
rlabel metal2 346948 556580 346948 556580 0 la_data_in[32]
rlabel via2 232070 518925 232070 518925 0 la_data_in[33]
rlabel metal2 232070 505223 232070 505223 0 la_data_in[34]
rlabel metal2 250010 1911 250010 1911 0 la_data_in[35]
rlabel metal2 253506 2608 253506 2608 0 la_data_in[36]
rlabel metal2 257094 2676 257094 2676 0 la_data_in[37]
rlabel via1 254702 556189 254702 556189 0 la_data_in[38]
rlabel metal2 232070 553843 232070 553843 0 la_data_in[39]
rlabel metal2 136482 2064 136482 2064 0 la_data_in[3]
rlabel metal2 229954 449123 229954 449123 0 la_data_in[40]
rlabel metal2 271025 340 271025 340 0 la_data_in[41]
rlabel metal2 274850 2744 274850 2744 0 la_data_in[42]
rlabel metal3 452080 409428 452080 409428 0 la_data_in[43]
rlabel metal3 234378 355708 234378 355708 0 la_data_in[44]
rlabel metal2 285193 340 285193 340 0 la_data_in[45]
rlabel metal2 289018 2200 289018 2200 0 la_data_in[46]
rlabel metal2 292606 161966 292606 161966 0 la_data_in[47]
rlabel metal2 296102 3220 296102 3220 0 la_data_in[48]
rlabel metal2 269668 556580 269668 556580 0 la_data_in[49]
rlabel metal2 140070 2574 140070 2574 0 la_data_in[4]
rlabel metal2 448346 556580 448346 556580 0 la_data_in[50]
rlabel metal2 232070 482273 232070 482273 0 la_data_in[51]
rlabel metal2 310270 3475 310270 3475 0 la_data_in[52]
rlabel metal2 313858 3560 313858 3560 0 la_data_in[53]
rlabel metal2 236226 338028 236226 338028 0 la_data_in[54]
rlabel metal2 320705 340 320705 340 0 la_data_in[55]
rlabel metal2 232070 501109 232070 501109 0 la_data_in[56]
rlabel metal2 328026 2115 328026 2115 0 la_data_in[57]
rlabel metal2 331469 340 331469 340 0 la_data_in[58]
rlabel metal2 334873 340 334873 340 0 la_data_in[59]
rlabel metal2 369488 556580 369488 556580 0 la_data_in[5]
rlabel metal2 409998 160475 409998 160475 0 la_data_in[60]
rlabel metal2 342194 1928 342194 1928 0 la_data_in[61]
rlabel metal2 345545 340 345545 340 0 la_data_in[62]
rlabel metal2 349232 16560 349232 16560 0 la_data_in[63]
rlabel metal2 352452 16560 352452 16560 0 la_data_in[64]
rlabel metal2 232070 484993 232070 484993 0 la_data_in[65]
rlabel metal2 464002 448324 464002 448324 0 la_data_in[66]
rlabel metal2 216614 231608 216614 231608 0 la_data_in[67]
rlabel metal3 233412 508028 233412 508028 0 la_data_in[68]
rlabel metal2 370385 340 370385 340 0 la_data_in[69]
rlabel metal3 452632 405348 452632 405348 0 la_data_in[6]
rlabel metal1 412850 333506 412850 333506 0 la_data_in[70]
rlabel metal3 452816 526388 452816 526388 0 la_data_in[71]
rlabel metal1 429548 559334 429548 559334 0 la_data_in[72]
rlabel metal2 384553 340 384553 340 0 la_data_in[73]
rlabel metal2 388049 340 388049 340 0 la_data_in[74]
rlabel metal2 391874 1911 391874 1911 0 la_data_in[75]
rlabel metal2 395048 16560 395048 16560 0 la_data_in[76]
rlabel metal1 438978 559402 438978 559402 0 la_data_in[77]
rlabel metal2 347898 160509 347898 160509 0 la_data_in[78]
rlabel metal2 405904 16560 405904 16560 0 la_data_in[79]
rlabel metal2 346548 338028 346548 338028 0 la_data_in[7]
rlabel metal3 233780 364548 233780 364548 0 la_data_in[80]
rlabel metal2 444406 160407 444406 160407 0 la_data_in[81]
rlabel metal2 463910 212432 463910 212432 0 la_data_in[82]
rlabel metal2 464094 448460 464094 448460 0 la_data_in[83]
rlabel metal2 423798 2268 423798 2268 0 la_data_in[84]
rlabel metal2 427294 2200 427294 2200 0 la_data_in[85]
rlabel metal2 430882 1911 430882 1911 0 la_data_in[86]
rlabel metal2 462438 281554 462438 281554 0 la_data_in[87]
rlabel metal2 463818 281248 463818 281248 0 la_data_in[88]
rlabel metal2 370944 556706 370944 556706 0 la_data_in[89]
rlabel metal2 154001 340 154001 340 0 la_data_in[8]
rlabel metal2 444498 16899 444498 16899 0 la_data_in[90]
rlabel metal3 234033 467228 234033 467228 0 la_data_in[91]
rlabel metal2 464278 420410 464278 420410 0 la_data_in[92]
rlabel metal2 332426 556580 332426 556580 0 la_data_in[93]
rlabel metal3 233941 437308 233941 437308 0 la_data_in[94]
rlabel metal2 462806 3627 462806 3627 0 la_data_in[95]
rlabel metal2 466065 340 466065 340 0 la_data_in[96]
rlabel metal2 387212 556580 387212 556580 0 la_data_in[97]
rlabel metal2 325726 169383 325726 169383 0 la_data_in[98]
rlabel metal3 233389 512108 233389 512108 0 la_data_in[99]
rlabel metal2 157596 16560 157596 16560 0 la_data_in[9]
rlabel metal2 366912 556580 366912 556580 0 la_data_out[0]
rlabel metal2 481758 1826 481758 1826 0 la_data_out[100]
rlabel metal2 485017 340 485017 340 0 la_data_out[101]
rlabel metal2 276200 338028 276200 338028 0 la_data_out[102]
rlabel metal3 452724 392428 452724 392428 0 la_data_out[103]
rlabel metal2 425852 556580 425852 556580 0 la_data_out[104]
rlabel metal3 452632 371348 452632 371348 0 la_data_out[105]
rlabel metal2 503010 3627 503010 3627 0 la_data_out[106]
rlabel metal2 489210 234260 489210 234260 0 la_data_out[107]
rlabel metal2 465750 245990 465750 245990 0 la_data_out[108]
rlabel metal2 513491 340 513491 340 0 la_data_out[109]
rlabel metal2 162281 340 162281 340 0 la_data_out[10]
rlabel metal3 233136 431868 233136 431868 0 la_data_out[110]
rlabel metal2 503010 196316 503010 196316 0 la_data_out[111]
rlabel metal3 233849 406708 233849 406708 0 la_data_out[112]
rlabel metal2 527528 16560 527528 16560 0 la_data_out[113]
rlabel metal2 253522 556580 253522 556580 0 la_data_out[114]
rlabel metal3 452632 369988 452632 369988 0 la_data_out[115]
rlabel metal2 538331 340 538331 340 0 la_data_out[116]
rlabel metal2 541512 16560 541512 16560 0 la_data_out[117]
rlabel metal2 545514 2268 545514 2268 0 la_data_out[118]
rlabel metal2 548865 340 548865 340 0 la_data_out[119]
rlabel metal2 463082 368934 463082 368934 0 la_data_out[11]
rlabel metal3 233757 388348 233757 388348 0 la_data_out[120]
rlabel metal1 438288 291822 438288 291822 0 la_data_out[121]
rlabel metal1 231380 346426 231380 346426 0 la_data_out[122]
rlabel metal2 563270 1962 563270 1962 0 la_data_out[123]
rlabel metal2 566352 16560 566352 16560 0 la_data_out[124]
rlabel metal1 405858 561714 405858 561714 0 la_data_out[125]
rlabel metal2 573705 340 573705 340 0 la_data_out[126]
rlabel metal2 577438 1860 577438 1860 0 la_data_out[127]
rlabel metal2 307970 168703 307970 168703 0 la_data_out[12]
rlabel metal2 172953 340 172953 340 0 la_data_out[13]
rlabel metal2 232070 545615 232070 545615 0 la_data_out[14]
rlabel metal2 179860 16560 179860 16560 0 la_data_out[15]
rlabel metal1 319010 327726 319010 327726 0 la_data_out[16]
rlabel metal2 465474 394519 465474 394519 0 la_data_out[17]
rlabel metal2 190663 340 190663 340 0 la_data_out[18]
rlabel metal2 194442 2064 194442 2064 0 la_data_out[19]
rlabel metal1 293986 333234 293986 333234 0 la_data_out[1]
rlabel metal2 197662 16560 197662 16560 0 la_data_out[20]
rlabel metal1 329498 333370 329498 333370 0 la_data_out[21]
rlabel via2 232070 520285 232070 520285 0 la_data_out[22]
rlabel metal1 330648 180098 330648 180098 0 la_data_out[23]
rlabel metal2 211961 340 211961 340 0 la_data_out[24]
rlabel metal2 215503 340 215503 340 0 la_data_out[25]
rlabel metal2 232070 465477 232070 465477 0 la_data_out[26]
rlabel metal2 222778 1758 222778 1758 0 la_data_out[27]
rlabel metal2 226366 1911 226366 1911 0 la_data_out[28]
rlabel metal2 229862 3424 229862 3424 0 la_data_out[29]
rlabel metal2 134182 3254 134182 3254 0 la_data_out[2]
rlabel metal2 233358 16560 233358 16560 0 la_data_out[30]
rlabel metal2 236801 340 236801 340 0 la_data_out[31]
rlabel metal3 234654 438668 234654 438668 0 la_data_out[32]
rlabel metal2 372018 556580 372018 556580 0 la_data_out[33]
rlabel metal2 247618 3526 247618 3526 0 la_data_out[34]
rlabel metal2 251206 163394 251206 163394 0 la_data_out[35]
rlabel metal2 254465 340 254465 340 0 la_data_out[36]
rlabel metal2 430760 338028 430760 338028 0 la_data_out[37]
rlabel metal1 449834 336702 449834 336702 0 la_data_out[38]
rlabel metal2 450570 169523 450570 169523 0 la_data_out[39]
rlabel metal2 137441 340 137441 340 0 la_data_out[3]
rlabel metal2 268633 340 268633 340 0 la_data_out[40]
rlabel metal3 234930 369988 234930 369988 0 la_data_out[41]
rlabel metal2 276046 3186 276046 3186 0 la_data_out[42]
rlabel metal3 234332 359108 234332 359108 0 la_data_out[43]
rlabel metal3 233964 450228 233964 450228 0 la_data_out[44]
rlabel metal2 286626 2710 286626 2710 0 la_data_out[45]
rlabel metal2 290214 2166 290214 2166 0 la_data_out[46]
rlabel metal2 293710 3152 293710 3152 0 la_data_out[47]
rlabel metal2 229862 445621 229862 445621 0 la_data_out[48]
rlabel metal2 224894 282557 224894 282557 0 la_data_out[49]
rlabel metal2 141036 16560 141036 16560 0 la_data_out[4]
rlabel metal3 233918 422348 233918 422348 0 la_data_out[50]
rlabel metal2 307970 2744 307970 2744 0 la_data_out[51]
rlabel metal1 231472 367098 231472 367098 0 la_data_out[52]
rlabel metal2 315054 1962 315054 1962 0 la_data_out[53]
rlabel metal3 233182 476748 233182 476748 0 la_data_out[54]
rlabel metal2 322138 3356 322138 3356 0 la_data_out[55]
rlabel metal2 325634 1928 325634 1928 0 la_data_out[56]
rlabel metal2 329222 1775 329222 1775 0 la_data_out[57]
rlabel metal2 332718 1163 332718 1163 0 la_data_out[58]
rlabel metal3 233274 448868 233274 448868 0 la_data_out[59]
rlabel metal2 353480 338028 353480 338028 0 la_data_out[5]
rlabel metal2 350766 338028 350766 338028 0 la_data_out[60]
rlabel metal2 343153 340 343153 340 0 la_data_out[61]
rlabel metal3 234424 380188 234424 380188 0 la_data_out[62]
rlabel metal2 350474 1928 350474 1928 0 la_data_out[63]
rlabel metal2 353825 340 353825 340 0 la_data_out[64]
rlabel metal2 408526 161257 408526 161257 0 la_data_out[65]
rlabel metal2 429426 338028 429426 338028 0 la_data_out[66]
rlabel metal2 364642 1911 364642 1911 0 la_data_out[67]
rlabel metal2 367993 340 367993 340 0 la_data_out[68]
rlabel metal2 371726 2064 371726 2064 0 la_data_out[69]
rlabel metal2 148113 340 148113 340 0 la_data_out[6]
rlabel metal2 392074 338028 392074 338028 0 la_data_out[70]
rlabel metal2 378665 340 378665 340 0 la_data_out[71]
rlabel metal3 233366 548828 233366 548828 0 la_data_out[72]
rlabel metal2 385986 3458 385986 3458 0 la_data_out[73]
rlabel metal2 389344 16560 389344 16560 0 la_data_out[74]
rlabel metal2 392833 340 392833 340 0 la_data_out[75]
rlabel metal2 292698 298413 292698 298413 0 la_data_out[76]
rlabel metal1 231426 374170 231426 374170 0 la_data_out[77]
rlabel metal2 345154 338028 345154 338028 0 la_data_out[78]
rlabel metal2 232070 372657 232070 372657 0 la_data_out[79]
rlabel metal2 151846 1911 151846 1911 0 la_data_out[7]
rlabel metal2 410826 1911 410826 1911 0 la_data_out[80]
rlabel via1 291226 556427 291226 556427 0 la_data_out[81]
rlabel metal3 233688 354348 233688 354348 0 la_data_out[82]
rlabel metal1 231058 532746 231058 532746 0 la_data_out[83]
rlabel metal3 234056 412148 234056 412148 0 la_data_out[84]
rlabel metal2 428214 16560 428214 16560 0 la_data_out[85]
rlabel metal2 432078 2608 432078 2608 0 la_data_out[86]
rlabel metal2 435337 340 435337 340 0 la_data_out[87]
rlabel metal3 233596 376788 233596 376788 0 la_data_out[88]
rlabel metal3 445901 334084 445901 334084 0 la_data_out[89]
rlabel metal2 155020 16560 155020 16560 0 la_data_out[8]
rlabel metal3 232653 527748 232653 527748 0 la_data_out[90]
rlabel metal2 449834 1792 449834 1792 0 la_data_out[91]
rlabel metal2 333592 556672 333592 556672 0 la_data_out[92]
rlabel metal3 233113 550188 233113 550188 0 la_data_out[93]
rlabel metal2 460039 340 460039 340 0 la_data_out[94]
rlabel metal2 464002 9476 464002 9476 0 la_data_out[95]
rlabel metal2 466992 16560 466992 16560 0 la_data_out[96]
rlabel metal2 470849 340 470849 340 0 la_data_out[97]
rlabel metal2 449680 556580 449680 556580 0 la_data_out[98]
rlabel metal1 231012 444414 231012 444414 0 la_data_out[99]
rlabel metal2 158838 16560 158838 16560 0 la_data_out[9]
rlabel metal2 405552 556580 405552 556580 0 la_oenb[0]
rlabel metal2 482625 340 482625 340 0 la_oenb[100]
rlabel metal2 486450 1962 486450 1962 0 la_oenb[101]
rlabel metal2 334098 181113 334098 181113 0 la_oenb[102]
rlabel metal2 493297 340 493297 340 0 la_oenb[103]
rlabel metal2 443240 556580 443240 556580 0 la_oenb[104]
rlabel metal2 500618 1962 500618 1962 0 la_oenb[105]
rlabel metal2 503969 340 503969 340 0 la_oenb[106]
rlabel metal2 291518 338028 291518 338028 0 la_oenb[107]
rlabel metal3 233090 389708 233090 389708 0 la_oenb[108]
rlabel metal1 395278 326774 395278 326774 0 la_oenb[109]
rlabel metal1 298310 557634 298310 557634 0 la_oenb[10]
rlabel metal3 232561 513468 232561 513468 0 la_oenb[110]
rlabel metal2 521771 340 521771 340 0 la_oenb[111]
rlabel metal2 525458 1911 525458 1911 0 la_oenb[112]
rlabel metal2 528809 340 528809 340 0 la_oenb[113]
rlabel metal2 500250 259250 500250 259250 0 la_oenb[114]
rlabel metal2 536130 2030 536130 2030 0 la_oenb[115]
rlabel metal2 539626 1996 539626 1996 0 la_oenb[116]
rlabel metal2 543214 4002 543214 4002 0 la_oenb[117]
rlabel metal2 546710 1928 546710 1928 0 la_oenb[118]
rlabel metal2 361606 300487 361606 300487 0 la_oenb[119]
rlabel metal1 346932 330446 346932 330446 0 la_oenb[11]
rlabel metal3 233826 435948 233826 435948 0 la_oenb[120]
rlabel metal2 525090 215798 525090 215798 0 la_oenb[121]
rlabel metal2 560641 340 560641 340 0 la_oenb[122]
rlabel metal2 564466 1894 564466 1894 0 la_oenb[123]
rlabel metal3 368989 557804 368989 557804 0 la_oenb[124]
rlabel metal2 313460 338028 313460 338028 0 la_oenb[125]
rlabel metal3 405674 559844 405674 559844 0 la_oenb[126]
rlabel metal3 232469 414868 232469 414868 0 la_oenb[127]
rlabel metal2 170561 340 170561 340 0 la_oenb[12]
rlabel metal2 174103 340 174103 340 0 la_oenb[13]
rlabel metal2 177882 4036 177882 4036 0 la_oenb[14]
rlabel metal2 181233 340 181233 340 0 la_oenb[15]
rlabel metal2 184966 5991 184966 5991 0 la_oenb[16]
rlabel metal1 272090 557974 272090 557974 0 la_oenb[17]
rlabel metal2 232070 390813 232070 390813 0 la_oenb[18]
rlabel metal2 195401 340 195401 340 0 la_oenb[19]
rlabel metal2 131790 3356 131790 3356 0 la_oenb[1]
rlabel metal2 198943 340 198943 340 0 la_oenb[20]
rlabel metal2 248538 160509 248538 160509 0 la_oenb[21]
rlabel metal2 206218 3492 206218 3492 0 la_oenb[22]
rlabel metal2 209806 3627 209806 3627 0 la_oenb[23]
rlabel metal2 212980 16560 212980 16560 0 la_oenb[24]
rlabel metal2 216798 16560 216798 16560 0 la_oenb[25]
rlabel metal2 220478 2710 220478 2710 0 la_oenb[26]
rlabel metal2 223783 340 223783 340 0 la_oenb[27]
rlabel metal2 385158 292905 385158 292905 0 la_oenb[28]
rlabel metal2 230782 16560 230782 16560 0 la_oenb[29]
rlabel metal2 135286 1911 135286 1911 0 la_oenb[2]
rlabel metal2 234646 23960 234646 23960 0 la_oenb[30]
rlabel metal2 237905 340 237905 340 0 la_oenb[31]
rlabel metal2 234646 335035 234646 335035 0 la_oenb[32]
rlabel metal3 233320 509388 233320 509388 0 la_oenb[33]
rlabel metal2 248623 340 248623 340 0 la_oenb[34]
rlabel metal2 232070 371297 232070 371297 0 la_oenb[35]
rlabel metal2 232070 443207 232070 443207 0 la_oenb[36]
rlabel metal1 356178 334730 356178 334730 0 la_oenb[37]
rlabel metal3 233734 403988 233734 403988 0 la_oenb[38]
rlabel metal4 235060 377808 235060 377808 0 la_oenb[39]
rlabel metal2 138874 2115 138874 2115 0 la_oenb[3]
rlabel metal2 269652 16560 269652 16560 0 la_oenb[40]
rlabel metal2 273509 340 273509 340 0 la_oenb[41]
rlabel metal2 276913 340 276913 340 0 la_oenb[42]
rlabel metal2 232070 452795 232070 452795 0 la_oenb[43]
rlabel metal1 369978 327794 369978 327794 0 la_oenb[44]
rlabel metal2 287585 340 287585 340 0 la_oenb[45]
rlabel metal3 233734 393788 233734 393788 0 la_oenb[46]
rlabel metal2 294492 16560 294492 16560 0 la_oenb[47]
rlabel metal3 234516 392428 234516 392428 0 la_oenb[48]
rlabel metal2 273486 338028 273486 338028 0 la_oenb[49]
rlabel metal2 293986 289437 293986 289437 0 la_oenb[4]
rlabel metal2 441738 161937 441738 161937 0 la_oenb[50]
rlabel metal2 309074 1622 309074 1622 0 la_oenb[51]
rlabel metal2 312425 340 312425 340 0 la_oenb[52]
rlabel metal3 234945 358428 234945 358428 0 la_oenb[53]
rlabel metal1 232760 349826 232760 349826 0 la_oenb[54]
rlabel metal2 232070 506583 232070 506583 0 la_oenb[55]
rlabel metal2 326593 340 326593 340 0 la_oenb[56]
rlabel metal2 330142 16560 330142 16560 0 la_oenb[57]
rlabel metal2 333914 1928 333914 1928 0 la_oenb[58]
rlabel metal2 337502 2183 337502 2183 0 la_oenb[59]
rlabel metal2 145721 340 145721 340 0 la_oenb[5]
rlabel metal3 452724 520948 452724 520948 0 la_oenb[60]
rlabel metal1 231472 382262 231472 382262 0 la_oenb[61]
rlabel metal2 348082 1911 348082 1911 0 la_oenb[62]
rlabel metal2 351670 2183 351670 2183 0 la_oenb[63]
rlabel metal2 460966 281588 460966 281588 0 la_oenb[64]
rlabel metal2 461426 448052 461426 448052 0 la_oenb[65]
rlabel metal2 232070 352461 232070 352461 0 la_oenb[66]
rlabel metal2 365838 3407 365838 3407 0 la_oenb[67]
rlabel metal2 369012 16560 369012 16560 0 la_oenb[68]
rlabel metal2 237560 338028 237560 338028 0 la_oenb[69]
rlabel metal2 405030 195840 405030 195840 0 la_oenb[6]
rlabel metal1 231426 374034 231426 374034 0 la_oenb[70]
rlabel metal2 379769 340 379769 340 0 la_oenb[71]
rlabel metal3 235060 491829 235060 491829 0 la_oenb[72]
rlabel metal1 230966 485826 230966 485826 0 la_oenb[73]
rlabel metal2 390632 16560 390632 16560 0 la_oenb[74]
rlabel metal1 230736 429182 230736 429182 0 la_oenb[75]
rlabel metal2 231978 415837 231978 415837 0 la_oenb[76]
rlabel metal2 232070 397681 232070 397681 0 la_oenb[77]
rlabel metal2 404846 2064 404846 2064 0 la_oenb[78]
rlabel metal2 408434 1860 408434 1860 0 la_oenb[79]
rlabel metal2 153042 2064 153042 2064 0 la_oenb[7]
rlabel metal2 232070 510697 232070 510697 0 la_oenb[80]
rlabel metal1 433596 334798 433596 334798 0 la_oenb[81]
rlabel metal2 462714 437376 462714 437376 0 la_oenb[82]
rlabel metal2 232070 462757 232070 462757 0 la_oenb[83]
rlabel metal2 232070 345627 232070 345627 0 la_oenb[84]
rlabel metal2 429449 340 429449 340 0 la_oenb[85]
rlabel metal2 433274 1724 433274 1724 0 la_oenb[86]
rlabel metal2 309550 556580 309550 556580 0 la_oenb[87]
rlabel metal2 440312 16560 440312 16560 0 la_oenb[88]
rlabel metal2 443854 2948 443854 2948 0 la_oenb[89]
rlabel metal2 156393 340 156393 340 0 la_oenb[8]
rlabel metal2 447304 16560 447304 16560 0 la_oenb[90]
rlabel metal2 450938 1758 450938 1758 0 la_oenb[91]
rlabel metal2 454526 3627 454526 3627 0 la_oenb[92]
rlabel metal3 235060 531609 235060 531609 0 la_oenb[93]
rlabel metal2 461610 1911 461610 1911 0 la_oenb[94]
rlabel metal1 464784 9622 464784 9622 0 la_oenb[95]
rlabel metal2 468457 340 468457 340 0 la_oenb[96]
rlabel metal3 452724 527748 452724 527748 0 la_oenb[97]
rlabel metal2 295366 203893 295366 203893 0 la_oenb[98]
rlabel metal3 452724 348908 452724 348908 0 la_oenb[99]
rlabel metal2 160126 275492 160126 275492 0 la_oenb[9]
rlabel metal4 235244 352512 235244 352512 0 user_irq[0]
rlabel metal3 235060 542897 235060 542897 0 user_irq[1]
rlabel metal2 583418 1843 583418 1843 0 user_irq[2]
rlabel metal2 361 340 361 340 0 wb_clk_i
rlabel metal2 1557 340 1557 340 0 wb_rst_i
rlabel metal2 2898 83307 2898 83307 0 wbs_ack_o
rlabel metal1 165646 561782 165646 561782 0 wbs_adr_i[0]
rlabel metal2 274820 556580 274820 556580 0 wbs_adr_i[10]
rlabel metal2 232070 502469 232070 502469 0 wbs_adr_i[11]
rlabel metal2 255346 294265 255346 294265 0 wbs_adr_i[12]
rlabel metal2 232070 464117 232070 464117 0 wbs_adr_i[13]
rlabel metal2 61817 340 61817 340 0 wbs_adr_i[14]
rlabel metal2 65313 340 65313 340 0 wbs_adr_i[15]
rlabel metal2 383794 338028 383794 338028 0 wbs_adr_i[16]
rlabel metal3 264385 315316 264385 315316 0 wbs_adr_i[17]
rlabel metal2 76077 340 76077 340 0 wbs_adr_i[18]
rlabel metal2 79481 340 79481 340 0 wbs_adr_i[19]
rlabel metal2 327122 556580 327122 556580 0 wbs_adr_i[1]
rlabel metal2 232070 410363 232070 410363 0 wbs_adr_i[20]
rlabel metal2 366114 336821 366114 336821 0 wbs_adr_i[21]
rlabel metal1 423338 336702 423338 336702 0 wbs_adr_i[22]
rlabel metal2 93978 8099 93978 8099 0 wbs_adr_i[23]
rlabel metal2 97060 16560 97060 16560 0 wbs_adr_i[24]
rlabel metal2 100917 340 100917 340 0 wbs_adr_i[25]
rlabel metal2 104321 340 104321 340 0 wbs_adr_i[26]
rlabel metal2 234738 555798 234738 555798 0 wbs_adr_i[27]
rlabel metal2 111642 1894 111642 1894 0 wbs_adr_i[28]
rlabel metal2 114993 340 114993 340 0 wbs_adr_i[29]
rlabel metal2 17066 1724 17066 1724 0 wbs_adr_i[2]
rlabel metal2 118818 3627 118818 3627 0 wbs_adr_i[30]
rlabel metal2 121900 16560 121900 16560 0 wbs_adr_i[31]
rlabel metal2 21850 1860 21850 1860 0 wbs_adr_i[3]
rlabel metal2 232806 547511 232806 547511 0 wbs_adr_i[4]
rlabel via2 232070 375411 232070 375411 0 wbs_adr_i[5]
rlabel metal2 306468 338028 306468 338028 0 wbs_adr_i[6]
rlabel metal2 36977 340 36977 340 0 wbs_adr_i[7]
rlabel metal2 40473 340 40473 340 0 wbs_adr_i[8]
rlabel metal2 44298 158515 44298 158515 0 wbs_adr_i[9]
rlabel metal2 3903 340 3903 340 0 wbs_cyc_i
rlabel metal4 235796 555628 235796 555628 0 wbs_dat_i[0]
rlabel metal2 232070 461363 232070 461363 0 wbs_dat_i[10]
rlabel metal2 232070 477819 232070 477819 0 wbs_dat_i[11]
rlabel metal2 55660 16560 55660 16560 0 wbs_dat_i[12]
rlabel metal2 59517 340 59517 340 0 wbs_dat_i[13]
rlabel metal2 62698 16560 62698 16560 0 wbs_dat_i[14]
rlabel metal2 66516 16560 66516 16560 0 wbs_dat_i[15]
rlabel metal2 232070 349707 232070 349707 0 wbs_dat_i[16]
rlabel metal1 289478 559266 289478 559266 0 wbs_dat_i[17]
rlabel metal2 77418 5328 77418 5328 0 wbs_dat_i[18]
rlabel metal2 80500 16560 80500 16560 0 wbs_dat_i[19]
rlabel metal2 21390 169898 21390 169898 0 wbs_dat_i[1]
rlabel metal2 84357 340 84357 340 0 wbs_dat_i[20]
rlabel metal2 234922 555985 234922 555985 0 wbs_dat_i[21]
rlabel metal2 232070 428485 232070 428485 0 wbs_dat_i[22]
rlabel metal2 94983 340 94983 340 0 wbs_dat_i[23]
rlabel metal2 98433 340 98433 340 0 wbs_dat_i[24]
rlabel metal2 102212 16560 102212 16560 0 wbs_dat_i[25]
rlabel metal2 232438 554166 232438 554166 0 wbs_dat_i[26]
rlabel metal2 217350 285600 217350 285600 0 wbs_dat_i[27]
rlabel metal2 112838 4104 112838 4104 0 wbs_dat_i[28]
rlabel metal2 116196 16560 116196 16560 0 wbs_dat_i[29]
rlabel metal2 18262 1894 18262 1894 0 wbs_dat_i[2]
rlabel metal2 119370 16560 119370 16560 0 wbs_dat_i[30]
rlabel via2 232070 423691 232070 423691 0 wbs_dat_i[31]
rlabel metal2 22809 340 22809 340 0 wbs_dat_i[3]
rlabel metal2 269330 183901 269330 183901 0 wbs_dat_i[4]
rlabel metal2 31089 340 31089 340 0 wbs_dat_i[5]
rlabel metal2 232070 338759 232070 338759 0 wbs_dat_i[6]
rlabel metal2 367034 558705 367034 558705 0 wbs_dat_i[7]
rlabel metal2 41676 16560 41676 16560 0 wbs_dat_i[8]
rlabel metal2 45303 340 45303 340 0 wbs_dat_i[9]
rlabel metal2 251298 303921 251298 303921 0 wbs_dat_o[0]
rlabel metal1 254196 312562 254196 312562 0 wbs_dat_o[10]
rlabel metal2 53774 2608 53774 2608 0 wbs_dat_o[11]
rlabel metal2 57033 340 57033 340 0 wbs_dat_o[12]
rlabel metal2 60858 3627 60858 3627 0 wbs_dat_o[13]
rlabel metal2 63940 16560 63940 16560 0 wbs_dat_o[14]
rlabel metal2 67797 340 67797 340 0 wbs_dat_o[15]
rlabel metal1 226458 235246 226458 235246 0 wbs_dat_o[16]
rlabel metal2 74796 16560 74796 16560 0 wbs_dat_o[17]
rlabel metal2 78423 340 78423 340 0 wbs_dat_o[18]
rlabel metal2 81873 340 81873 340 0 wbs_dat_o[19]
rlabel metal2 405858 274953 405858 274953 0 wbs_dat_o[1]
rlabel via2 232070 426445 232070 426445 0 wbs_dat_o[20]
rlabel via2 232070 516171 232070 516171 0 wbs_dat_o[21]
rlabel metal2 92637 340 92637 340 0 wbs_dat_o[22]
rlabel metal2 96041 340 96041 340 0 wbs_dat_o[23]
rlabel metal2 99636 16560 99636 16560 0 wbs_dat_o[24]
rlabel metal2 103362 2030 103362 2030 0 wbs_dat_o[25]
rlabel metal2 106713 340 106713 340 0 wbs_dat_o[26]
rlabel metal2 292208 556580 292208 556580 0 wbs_dat_o[27]
rlabel metal2 114034 1996 114034 1996 0 wbs_dat_o[28]
rlabel metal2 117477 340 117477 340 0 wbs_dat_o[29]
rlabel metal2 19412 16560 19412 16560 0 wbs_dat_o[2]
rlabel metal2 120881 340 120881 340 0 wbs_dat_o[30]
rlabel metal4 463772 422076 463772 422076 0 wbs_dat_o[31]
rlabel metal2 24242 1962 24242 1962 0 wbs_dat_o[3]
rlabel metal2 28934 1928 28934 1928 0 wbs_dat_o[4]
rlabel metal2 32430 1911 32430 1911 0 wbs_dat_o[5]
rlabel metal2 36018 3627 36018 3627 0 wbs_dat_o[6]
rlabel metal2 39606 1979 39606 1979 0 wbs_dat_o[7]
rlabel metal2 42957 340 42957 340 0 wbs_dat_o[8]
rlabel metal2 373352 556580 373352 556580 0 wbs_dat_o[9]
rlabel metal2 232070 541501 232070 541501 0 wbs_sel_i[0]
rlabel metal1 137356 557770 137356 557770 0 wbs_sel_i[1]
rlabel metal2 20654 1843 20654 1843 0 wbs_sel_i[2]
rlabel metal2 232070 385339 232070 385339 0 wbs_sel_i[3]
rlabel metal2 232070 521985 232070 521985 0 wbs_stb_i
rlabel metal2 6249 340 6249 340 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
