##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Sun Jun  5 21:30:06 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO soc_now_caravel_top
  CLASS BLOCK ;
  SIZE 1200.140000 BY 930.580000 ;
  FOREIGN soc_now_caravel_top 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9573 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.6255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 80.164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 428.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.4482 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.556 LAYER met4  ;
    ANTENNAMAXAREACAR 77.6376 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 419.405 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.248122 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 2.330000 0.000000 2.470000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.9764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 170.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.708 LAYER met3  ;
    ANTENNAMAXAREACAR 111.102 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 564.925 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.403446 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 0.530000 0.800000 0.830000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.330000 0.000000 251.470000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.530000 0.000000 84.670000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.730000 0.000000 253.870000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.830000 0.000000 248.970000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.430000 0.000000 246.570000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.130000 0.000000 244.270000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.630000 0.000000 241.770000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.830000 0.000000 161.970000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.430000 0.000000 159.570000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.030000 0.000000 157.170000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.630000 0.000000 154.770000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.130000 0.000000 152.270000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.730000 0.000000 149.870000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.330000 0.000000 147.470000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.930000 0.000000 145.070000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.530000 0.000000 142.670000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.030000 0.000000 140.170000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630000 0.000000 137.770000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.230000 0.000000 135.370000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.830000 0.000000 132.970000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.430000 0.000000 130.570000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.930000 0.000000 128.070000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.530000 0.000000 125.670000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.230000 0.000000 123.370000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.730000 0.000000 120.870000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.330000 0.000000 118.470000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.930000 0.000000 116.070000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.530000 0.000000 113.670000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.130000 0.000000 111.270000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.630000 0.000000 108.770000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.230000 0.000000 106.370000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.830000 0.000000 103.970000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.430000 0.000000 101.570000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.030000 0.000000 99.170000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.630000 0.000000 96.770000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.130000 0.000000 94.270000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.730000 0.000000 91.870000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330000 0.000000 89.470000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.930000 0.000000 87.070000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.030000 0.000000 82.170000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.630000 0.000000 79.770000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230000 0.000000 77.370000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.830000 0.000000 74.970000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.430000 0.000000 72.570000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.930000 0.000000 70.070000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.530000 0.000000 67.670000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.130000 0.000000 65.270000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.730000 0.000000 62.870000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.330000 0.000000 60.470000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.830000 0.000000 57.970000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.430000 0.000000 55.570000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.030000 0.000000 53.170000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.630000 0.000000 50.770000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.230000 0.000000 48.370000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.830000 0.000000 45.970000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330000 0.000000 43.470000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.930000 0.000000 41.070000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.530000 0.000000 38.670000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.130000 0.000000 36.270000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.730000 0.000000 33.870000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.230000 0.000000 31.370000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.830000 0.000000 28.970000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.430000 0.000000 26.570000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.030000 0.000000 24.170000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.630000 0.000000 21.770000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.130000 0.000000 19.270000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.730000 0.000000 16.870000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.330000 0.000000 14.470000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.930000 0.000000 12.070000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.530000 0.000000 9.670000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.130000 0.000000 7.270000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 4.630000 0.000000 4.770000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.230000 0.000000 239.370000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 236.830000 0.000000 236.970000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 234.430000 0.000000 234.570000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 232.030000 0.000000 232.170000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.530000 0.000000 229.670000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 227.130000 0.000000 227.270000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 224.730000 0.000000 224.870000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 222.330000 0.000000 222.470000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 219.930000 0.000000 220.070000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 217.430000 0.000000 217.570000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 215.030000 0.000000 215.170000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 212.630000 0.000000 212.770000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 210.230000 0.000000 210.370000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 207.830000 0.000000 207.970000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 205.330000 0.000000 205.470000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 202.930000 0.000000 203.070000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 200.530000 0.000000 200.670000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 198.130000 0.000000 198.270000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 195.730000 0.000000 195.870000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 193.330000 0.000000 193.470000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.830000 0.000000 190.970000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 188.430000 0.000000 188.570000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.030000 0.000000 186.170000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 183.630000 0.000000 183.770000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 181.230000 0.000000 181.370000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 178.730000 0.000000 178.870000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 176.330000 0.000000 176.470000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 173.930000 0.000000 174.070000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 171.530000 0.000000 171.670000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 169.130000 0.000000 169.270000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.630000 0.000000 166.770000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 164.230000 0.000000 164.370000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.230000 0.000000 563.370000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830000 0.000000 560.970000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.330000 0.000000 558.470000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.930000 0.000000 556.070000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.530000 0.000000 553.670000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.130000 0.000000 551.270000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.730000 0.000000 548.870000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.330000 0.000000 546.470000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.830000 0.000000 543.970000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.430000 0.000000 541.570000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.030000 0.000000 539.170000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.630000 0.000000 536.770000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.230000 0.000000 534.370000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.730000 0.000000 531.870000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.330000 0.000000 529.470000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.930000 0.000000 527.070000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.530000 0.000000 524.670000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.130000 0.000000 522.270000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.630000 0.000000 519.770000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.230000 0.000000 517.370000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830000 0.000000 514.970000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.430000 0.000000 512.570000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.030000 0.000000 510.170000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.530000 0.000000 507.670000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.130000 0.000000 505.270000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.730000 0.000000 502.870000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.330000 0.000000 500.470000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.930000 0.000000 498.070000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.530000 0.000000 495.670000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.030000 0.000000 493.170000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.630000 0.000000 490.770000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.230000 0.000000 488.370000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.830000 0.000000 485.970000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.430000 0.000000 483.570000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.030000 0.000000 481.170000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.630000 0.000000 478.770000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.230000 0.000000 476.370000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.730000 0.000000 473.870000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.330000 0.000000 471.470000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.930000 0.000000 469.070000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530000 0.000000 466.670000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.130000 0.000000 464.270000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.630000 0.000000 461.770000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.230000 0.000000 459.370000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.830000 0.000000 456.970000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.430000 0.000000 454.570000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.030000 0.000000 452.170000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.630000 0.000000 449.770000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.130000 0.000000 447.270000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.730000 0.000000 444.870000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.330000 0.000000 442.470000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.930000 0.000000 440.070000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.530000 0.000000 437.670000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.030000 0.000000 435.170000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.630000 0.000000 432.770000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.230000 0.000000 430.370000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.830000 0.000000 427.970000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.430000 0.000000 425.570000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.930000 0.000000 423.070000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530000 0.000000 420.670000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.130000 0.000000 418.270000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.730000 0.000000 415.870000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.330000 0.000000 413.470000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.830000 0.000000 410.970000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.430000 0.000000 408.570000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.030000 0.000000 406.170000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.630000 0.000000 403.770000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.230000 0.000000 401.370000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.830000 0.000000 398.970000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.330000 0.000000 396.470000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.930000 0.000000 394.070000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.530000 0.000000 391.670000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.130000 0.000000 389.270000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.730000 0.000000 386.870000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.230000 0.000000 384.370000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.830000 0.000000 381.970000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.430000 0.000000 379.570000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.030000 0.000000 377.170000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.630000 0.000000 374.770000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.130000 0.000000 372.270000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.730000 0.000000 369.870000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.330000 0.000000 367.470000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.930000 0.000000 365.070000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.530000 0.000000 362.670000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.130000 0.000000 360.270000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.730000 0.000000 357.870000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.330000 0.000000 355.470000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.830000 0.000000 352.970000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.430000 0.000000 350.570000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.030000 0.000000 348.170000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.630000 0.000000 345.770000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.230000 0.000000 343.370000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.830000 0.000000 340.970000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.330000 0.000000 338.470000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.930000 0.000000 336.070000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.530000 0.000000 333.670000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.130000 0.000000 331.270000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.730000 0.000000 328.870000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230000 0.000000 326.370000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.830000 0.000000 323.970000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.430000 0.000000 321.570000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.030000 0.000000 319.170000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.630000 0.000000 316.770000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.130000 0.000000 314.270000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.730000 0.000000 311.870000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.330000 0.000000 309.470000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.930000 0.000000 307.070000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.530000 0.000000 304.670000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.130000 0.000000 302.270000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.630000 0.000000 299.770000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.230000 0.000000 297.370000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.830000 0.000000 294.970000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.942 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.2262 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 292.430000 0.000000 292.570000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1124 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.9722 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 290.030000 0.000000 290.170000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.521 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 16.248 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.8095 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 287.530000 0.000000 287.670000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1073 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.9203 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 285.130000 0.000000 285.270000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 9.23495 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.0556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 282.730000 0.000000 282.870000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0748 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.148 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 10.9112 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.1232 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 280.330000 0.000000 280.470000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7884 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.834 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.83232 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.9788 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 277.930000 0.000000 278.070000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.264 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.38929 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.7354 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 275.430000 0.000000 275.570000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0662 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.115 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 4.89716 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.7075 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.289606 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 273.030000 0.000000 273.170000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1642 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.66667 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.2727 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 270.630000 0.000000 270.770000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 5.42494 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.0912 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 268.230000 0.000000 268.370000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 7.82606 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.0697 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 265.830000 0.000000 265.970000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.194 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 6.97883 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.7251 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 263.330000 0.000000 263.470000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3104 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.326 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 8.2295 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 260.930000 0.000000 261.070000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8206 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.995 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.38633 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.301 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.147071 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 258.530000 0.000000 258.670000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.412 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 6.1017 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.1372 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 256.130000 0.000000 256.270000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.984 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.115 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.104 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.488 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 555.644 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 872.630000 0.000000 872.770000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.0855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.1649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.621 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 556.16 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 870.230000 0.000000 870.370000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.0855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.1649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.621 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 556.16 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 867.830000 0.000000 867.970000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.0855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.1649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.621 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 556.16 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 865.430000 0.000000 865.570000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.0855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.1649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.621 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 556.16 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 863.030000 0.000000 863.170000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.0855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.1649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.621 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 556.16 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 860.530000 0.000000 860.670000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.0855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.1649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.621 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 556.16 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 858.130000 0.000000 858.270000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.033 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.1649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.354 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 555.893 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 855.730000 0.000000 855.870000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.033 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.1649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.354 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 555.893 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 853.330000 0.000000 853.470000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.0855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.1649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.621 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 556.16 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 850.930000 0.000000 851.070000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.0855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 50.6641 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 249.328 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 105.037 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 565.868 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 848.530000 0.000000 848.670000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.1065 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.2397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.728 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.612 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 556.267 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 846.130000 0.000000 846.270000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 843.730000 0.000000 843.870000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 841.330000 0.000000 841.470000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 838.830000 0.000000 838.970000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 836.430000 0.000000 836.570000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 123.711 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 611.082 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.241315 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 834.030000 0.000000 834.170000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 831.630000 0.000000 831.770000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 829.230000 0.000000 829.370000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 826.730000 0.000000 826.870000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 824.330000 0.000000 824.470000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 821.930000 0.000000 822.070000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 819.530000 0.000000 819.670000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 817.130000 0.000000 817.270000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 814.630000 0.000000 814.770000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 812.230000 0.000000 812.370000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 809.830000 0.000000 809.970000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 807.430000 0.000000 807.570000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 805.030000 0.000000 805.170000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 802.530000 0.000000 802.670000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 800.130000 0.000000 800.270000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 797.730000 0.000000 797.870000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 795.330000 0.000000 795.470000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 792.930000 0.000000 793.070000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 790.530000 0.000000 790.670000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 788.030000 0.000000 788.170000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 785.630000 0.000000 785.770000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 783.230000 0.000000 783.370000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 780.830000 0.000000 780.970000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 778.430000 0.000000 778.570000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 775.930000 0.000000 776.070000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 773.530000 0.000000 773.670000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 771.130000 0.000000 771.270000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 768.730000 0.000000 768.870000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 766.330000 0.000000 766.470000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 763.830000 0.000000 763.970000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 761.430000 0.000000 761.570000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 759.030000 0.000000 759.170000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 756.630000 0.000000 756.770000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 754.230000 0.000000 754.370000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.546 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.262 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 608.195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 751.730000 0.000000 751.870000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 749.330000 0.000000 749.470000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 746.930000 0.000000 747.070000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 744.530000 0.000000 744.670000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 742.130000 0.000000 742.270000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 739.730000 0.000000 739.870000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 737.230000 0.000000 737.370000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 734.830000 0.000000 734.970000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 732.430000 0.000000 732.570000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 730.030000 0.000000 730.170000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 727.630000 0.000000 727.770000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 725.230000 0.000000 725.370000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 722.830000 0.000000 722.970000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 720.430000 0.000000 720.570000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 717.930000 0.000000 718.070000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 715.530000 0.000000 715.670000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 713.130000 0.000000 713.270000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 710.730000 0.000000 710.870000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 708.330000 0.000000 708.470000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 705.830000 0.000000 705.970000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 703.430000 0.000000 703.570000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 701.030000 0.000000 701.170000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 698.630000 0.000000 698.770000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 696.230000 0.000000 696.370000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 693.830000 0.000000 693.970000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 691.330000 0.000000 691.470000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 688.930000 0.000000 689.070000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 686.530000 0.000000 686.670000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 684.130000 0.000000 684.270000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 681.730000 0.000000 681.870000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.62 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 679.230000 0.000000 679.370000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 676.830000 0.000000 676.970000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 674.430000 0.000000 674.570000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 672.030000 0.000000 672.170000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.205 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 669.630000 0.000000 669.770000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.0198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.374 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met2  ;
    ANTENNAMAXAREACAR 122.159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 607.39 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 667.130000 0.000000 667.270000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 664.730000 0.000000 664.870000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 662.330000 0.000000 662.470000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 659.930000 0.000000 660.070000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 657.530000 0.000000 657.670000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 655.030000 0.000000 655.170000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 652.630000 0.000000 652.770000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 650.230000 0.000000 650.370000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 647.830000 0.000000 647.970000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 645.430000 0.000000 645.570000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 643.030000 0.000000 643.170000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 640.530000 0.000000 640.670000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 638.130000 0.000000 638.270000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 635.730000 0.000000 635.870000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 633.330000 0.000000 633.470000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 630.930000 0.000000 631.070000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 628.430000 0.000000 628.570000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 626.030000 0.000000 626.170000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 623.630000 0.000000 623.770000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 621.230000 0.000000 621.370000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 618.830000 0.000000 618.970000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 616.330000 0.000000 616.470000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 613.930000 0.000000 614.070000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 611.530000 0.000000 611.670000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 609.130000 0.000000 609.270000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 606.730000 0.000000 606.870000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 604.330000 0.000000 604.470000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 601.930000 0.000000 602.070000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 599.530000 0.000000 599.670000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 597.130000 0.000000 597.270000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 594.630000 0.000000 594.770000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 592.230000 0.000000 592.370000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 589.830000 0.000000 589.970000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 587.430000 0.000000 587.570000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 585.030000 0.000000 585.170000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 582.530000 0.000000 582.670000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 580.130000 0.000000 580.270000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 577.730000 0.000000 577.870000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 575.330000 0.000000 575.470000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 572.930000 0.000000 573.070000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 570.430000 0.000000 570.570000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 568.030000 0.000000 568.170000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.2584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 565.630000 0.000000 565.770000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.230000 0.000000 1182.370000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.730000 0.000000 1179.870000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.330000 0.000000 1177.470000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.930000 0.000000 1175.070000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.530000 0.000000 1172.670000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.130000 0.000000 1170.270000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.630000 0.000000 1167.770000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.230000 0.000000 1165.370000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.830000 0.000000 1162.970000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.430000 0.000000 1160.570000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.030000 0.000000 1158.170000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.530000 0.000000 1155.670000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.130000 0.000000 1153.270000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.730000 0.000000 1150.870000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.330000 0.000000 1148.470000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.930000 0.000000 1146.070000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.430000 0.000000 1143.570000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.030000 0.000000 1141.170000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.630000 0.000000 1138.770000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.230000 0.000000 1136.370000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.830000 0.000000 1133.970000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.430000 0.000000 1131.570000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.930000 0.000000 1129.070000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.530000 0.000000 1126.670000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.130000 0.000000 1124.270000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.730000 0.000000 1121.870000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.330000 0.000000 1119.470000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.830000 0.000000 1116.970000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.430000 0.000000 1114.570000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.030000 0.000000 1112.170000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.630000 0.000000 1109.770000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.230000 0.000000 1107.370000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.730000 0.000000 1104.870000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.330000 0.000000 1102.470000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.930000 0.000000 1100.070000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.530000 0.000000 1097.670000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.130000 0.000000 1095.270000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.730000 0.000000 1092.870000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.330000 0.000000 1090.470000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.930000 0.000000 1088.070000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.530000 0.000000 1085.670000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.030000 0.000000 1083.170000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630000 0.000000 1080.770000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.230000 0.000000 1078.370000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.830000 0.000000 1075.970000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.430000 0.000000 1073.570000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.930000 0.000000 1071.070000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.530000 0.000000 1068.670000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.130000 0.000000 1066.270000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.730000 0.000000 1063.870000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.330000 0.000000 1061.470000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.830000 0.000000 1058.970000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.430000 0.000000 1056.570000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.030000 0.000000 1054.170000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.630000 0.000000 1051.770000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.230000 0.000000 1049.370000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.730000 0.000000 1046.870000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.330000 0.000000 1044.470000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.930000 0.000000 1042.070000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.530000 0.000000 1039.670000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.130000 0.000000 1037.270000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.730000 0.000000 1034.870000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.230000 0.000000 1032.370000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.830000 0.000000 1029.970000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.430000 0.000000 1027.570000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.030000 0.000000 1025.170000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.630000 0.000000 1022.770000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.130000 0.000000 1020.270000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.730000 0.000000 1017.870000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.330000 0.000000 1015.470000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.930000 0.000000 1013.070000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.530000 0.000000 1010.670000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.030000 0.000000 1008.170000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.630000 0.000000 1005.770000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.230000 0.000000 1003.370000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.830000 0.000000 1000.970000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.430000 0.000000 998.570000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.930000 0.000000 996.070000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.530000 0.000000 993.670000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.130000 0.000000 991.270000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.730000 0.000000 988.870000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330000 0.000000 986.470000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.930000 0.000000 984.070000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.430000 0.000000 981.570000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.030000 0.000000 979.170000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.630000 0.000000 976.770000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.230000 0.000000 974.370000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.830000 0.000000 971.970000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.430000 0.000000 969.570000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.030000 0.000000 967.170000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.630000 0.000000 964.770000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.130000 0.000000 962.270000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.730000 0.000000 959.870000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.330000 0.000000 957.470000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.930000 0.000000 955.070000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.530000 0.000000 952.670000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.030000 0.000000 950.170000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.630000 0.000000 947.770000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.230000 0.000000 945.370000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.830000 0.000000 942.970000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.430000 0.000000 940.570000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030000 0.000000 938.170000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.530000 0.000000 935.670000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.130000 0.000000 933.270000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.730000 0.000000 930.870000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.330000 0.000000 928.470000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.930000 0.000000 926.070000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.430000 0.000000 923.570000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.030000 0.000000 921.170000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.630000 0.000000 918.770000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.230000 0.000000 916.370000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.830000 0.000000 913.970000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.330000 0.000000 911.470000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.930000 0.000000 909.070000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.530000 0.000000 906.670000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.130000 0.000000 904.270000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.730000 0.000000 901.870000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.230000 0.000000 899.370000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.830000 0.000000 896.970000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.430000 0.000000 894.570000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030000 0.000000 892.170000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.630000 0.000000 889.770000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.230000 0.000000 887.370000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.730000 0.000000 884.870000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.330000 0.000000 882.470000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.930000 0.000000 880.070000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.530000 0.000000 877.670000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.130000 0.000000 875.270000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.0114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 75.5628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 403.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 145.577 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 702.642 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.782377 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.080000 0.800000 34.380000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.9594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 170.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.5377 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 414 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 149.214 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 786.058 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 85.320000 0.800000 85.620000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 180.936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 965.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.1246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 94.0067 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 499.374 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 136.560000 0.800000 136.860000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 100.862 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 537.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.4104 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 63.7372 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.101 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 204.880000 0.800000 205.180000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 121.601 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 648.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.2026 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 87.8879 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 463.269 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 273.200000 0.800000 273.500000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 240.242 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1281.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.3188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 45.3472 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 234.411 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.621614 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 341.520000 0.800000 341.820000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.1784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 300.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.8336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 123.339 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 645.412 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 409.840000 0.800000 410.140000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 159.393 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 850.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.9336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 96.9516 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 504.962 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 478.160000 0.800000 478.460000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 133.658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 713.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.0704 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 46.6847 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 245.965 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.782377 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 546.480000 0.800000 546.780000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 55.6823 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 270.127 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.675745 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 614.800000 0.800000 615.100000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 108.774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 580.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 26.9379 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 131.436 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 683.120000 0.800000 683.420000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.464 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 40.5297 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 200.644 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.464917 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 751.440000 0.800000 751.740000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 55.1972 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 277.596 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.643488 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 819.760000 0.800000 820.060000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.0094 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 57.6759 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.546 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 887.470000 0.800000 887.770000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.4837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 227.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 70.0086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 374.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 162.456 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 792.379 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.751262 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 67.930000 930.090000 68.070000 930.580000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 213.297 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met2  ;
    ANTENNAMAXAREACAR 67.2074 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 332.56 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 204.230000 930.090000 204.370000 930.580000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.6249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 212.846 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 88.6746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 473.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 194.721 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 991.36 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732726 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 340.430000 930.090000 340.570000 930.580000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.4187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 356.814 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.806 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.2088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 225.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 78.7461 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.384 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 476.630000 930.090000 476.770000 930.580000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 61.1975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 305.827 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.7334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 330.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 108.308 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 514.121 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 612.930000 930.090000 613.070000 930.580000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 70.2091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.767 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.3716 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 101.551 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 536.498 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 749.130000 930.090000 749.270000 930.580000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.6202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 172.403 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met2  ;
    ANTENNAMAXAREACAR 64.1745 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 314.398 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.497222 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 885.330000 930.090000 885.470000 930.580000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.2522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 155.337 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met2  ;
    ANTENNAMAXAREACAR 72.9367 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 353.952 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1021.530000 930.090000 1021.670000 930.580000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.4333 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 212.006 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 89.6357 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 445.639 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.879039 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1157.730000 930.090000 1157.870000 930.580000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7293 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.9728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 48.537 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.971 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.960948 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 869.170000 1200.140000 869.470000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 105.979 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 516.676 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.643488 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 799.630000 1200.140000 799.930000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 81.772 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 406.41 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.643488 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 730.090000 1200.140000 730.390000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 81.8092 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 408.215 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.643488 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 660.550000 1200.140000 660.850000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 54.6073 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 270.171 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.643488 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 591.010000 1200.140000 591.310000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.4294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 71.7107 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 357.286 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.643488 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 521.470000 1200.140000 521.770000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 37.93 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 189.816 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.464917 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 451.930000 1200.140000 452.230000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 86.7646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 462.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 36.5134 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 172.15 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 382.390000 1200.140000 382.690000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 116.274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 620.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 17.5219 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 84.333 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 312.850000 1200.140000 313.150000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 183.296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 977.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.0904 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 44.5279 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.829 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 260.390000 1200.140000 260.690000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 208.540000 1200.140000 208.840000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 156.080000 1200.140000 156.380000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 103.620000 1200.140000 103.920000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 51.770000 1200.140000 52.070000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.760000 0.000000 1200.060000 0.800000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.2954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 220.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 72.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 387.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 104.968 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 547.753 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 17.000000 0.800000 17.300000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.9524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.6108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 419.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 100.584 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 528.981 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 68.240000 0.800000 68.540000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.5428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 462.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 111.574 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 585.636 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.480000 0.800000 119.780000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 91.1566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 486.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.7536 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.96 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 187.800000 0.800000 188.100000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 152.993 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 815.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.4128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.672 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 256.120000 0.800000 256.420000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 115.67 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 616.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 324.440000 0.800000 324.740000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 118.535 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 632.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.2216 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.456 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 392.760000 0.800000 393.060000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.6144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 233.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.1658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 67.8041 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 350.115 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.470303 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 461.080000 0.800000 461.380000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 83.5654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 446.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.4754 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 109.145 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 574.991 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.470303 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 529.400000 0.800000 529.700000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 88.528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 474.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 206.25 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1087.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.450101 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 206.924 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1091.83 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.450101 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 597.720000 0.800000 598.020000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.9194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 60.9999 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 310.919 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.496162 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 666.040000 0.800000 666.340000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.4014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 83.9656 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 419.289 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.33899 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 734.360000 0.800000 734.660000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7583 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.4946 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 64.3327 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 339.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 802.070000 0.800000 802.370000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.4256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 143.126 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 763.107 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.450101 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 871.000000 0.800000 871.300000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.4352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 116.704 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 50.8287 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 249.269 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 33.930000 930.090000 34.070000 930.580000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.5007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.2245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.8844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 150.028 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 792.629 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.712727 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 170.130000 930.090000 170.270000 930.580000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.4184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.866 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 306.430000 930.090000 306.570000 930.580000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 72.3328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 361.438 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 442.630000 930.090000 442.770000 930.580000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 70.1069 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.87 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.5888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.944 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 578.830000 930.090000 578.970000 930.580000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.1375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.209 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 172.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 146.782 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 783.776 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 715.030000 930.090000 715.170000 930.580000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.4435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.521 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 189.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.0198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.0292 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 394.119 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423165 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 851.230000 930.090000 851.370000 930.580000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 85.3078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 426.195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 987.530000 930.090000 987.670000 930.580000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 83.5622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 417.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1123.730000 930.090000 1123.870000 930.580000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 886.860000 1200.140000 887.160000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.5564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 817.320000 1200.140000 817.620000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 747.780000 1200.140000 748.080000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.0744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 144.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 678.240000 1200.140000 678.540000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.8434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 608.700000 1200.140000 609.000000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.9814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.896 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 538.550000 1200.140000 538.850000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 469.010000 1200.140000 469.310000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 110.51 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 589.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 166.905 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 878.828 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352458 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 399.470000 1200.140000 399.770000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 117.275 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 625.464 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 172.617 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 912.532 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.443367 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 329.930000 1200.140000 330.230000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.7618 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 313.282 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 278.080000 1200.140000 278.380000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.3802 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.247 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 225.620000 1200.140000 225.920000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.3802 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.247 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 173.160000 1200.140000 173.460000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.3802 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.247 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 121.310000 1200.140000 121.610000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.7618 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 313.282 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 68.850000 1200.140000 69.150000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.7618 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 313.282 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 17.000000 1200.140000 17.300000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 71.0934 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 379.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1.250000 0.000000 1.550000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 51.160000 0.800000 51.460000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 102.400000 0.800000 102.700000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 60.1014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 320.536 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 170.720000 0.800000 171.020000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 60.6534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 323.48 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 239.040000 0.800000 239.340000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 307.360000 0.800000 307.660000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 49.8894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 266.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 375.680000 0.800000 375.980000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 444.000000 0.800000 444.300000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 512.320000 0.800000 512.620000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.9024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 580.640000 0.800000 580.940000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 66.0612 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 352.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 648.960000 0.800000 649.260000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.44 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 717.280000 0.800000 717.580000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 785.600000 0.800000 785.900000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3934 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.9068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 458.64 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 853.920000 0.800000 854.220000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 73.9316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 369.432 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1.030000 930.090000 1.170000 930.580000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 73.5422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 367.367 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 136.030000 930.090000 136.170000 930.580000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.7834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.691 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 272.330000 930.090000 272.470000 930.580000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.7684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.498 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 408.530000 930.090000 408.670000 930.580000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.1392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.588 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 544.730000 930.090000 544.870000 930.580000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.397 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.877 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 680.930000 930.090000 681.070000 930.580000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.141 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 817.230000 930.090000 817.370000 930.580000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.764 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 953.430000 930.090000 953.570000 930.580000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.554 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1089.630000 930.090000 1089.770000 930.580000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.0484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 903.940000 1200.140000 904.240000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.2914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 834.400000 1200.140000 834.700000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.0044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 764.860000 1200.140000 765.160000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.7644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 695.320000 1200.140000 695.620000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.7734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 132.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 625.780000 1200.140000 626.080000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 556.240000 1200.140000 556.540000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 486.700000 1200.140000 487.000000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 63.7824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 340.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 417.160000 1200.140000 417.460000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 347.620000 1200.140000 347.920000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 295.160000 1200.140000 295.460000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.3802 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.247 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 243.310000 1200.140000 243.610000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.3802 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.247 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 190.850000 1200.140000 191.150000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.3802 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.247 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 138.390000 1200.140000 138.690000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.7618 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 313.282 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 86.540000 1200.140000 86.840000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 53.7618 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 313.282 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 34.080000 1200.140000 34.380000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 153.640000 0.800000 153.940000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 221.960000 0.800000 222.260000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 290.280000 0.800000 290.580000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 358.600000 0.800000 358.900000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 426.920000 0.800000 427.220000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 495.240000 0.800000 495.540000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 563.560000 0.800000 563.860000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 631.880000 0.800000 632.180000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 700.200000 0.800000 700.500000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 768.520000 0.800000 768.820000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 836.840000 0.800000 837.140000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 904.550000 0.800000 904.850000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.030000 930.090000 102.170000 930.580000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.230000 930.090000 238.370000 930.580000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.430000 930.090000 374.570000 930.580000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.730000 930.090000 510.870000 930.580000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.930000 930.090000 647.070000 930.580000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.130000 930.090000 783.270000 930.580000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.430000 930.090000 919.570000 930.580000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.630000 930.090000 1055.770000 930.580000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.930000 930.090000 1191.070000 930.580000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 852.090000 1200.140000 852.390000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 782.550000 1200.140000 782.850000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 713.010000 1200.140000 713.310000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 643.470000 1200.140000 643.770000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 573.930000 1200.140000 574.230000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 503.780000 1200.140000 504.080000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 434.240000 1200.140000 434.540000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.340000 364.700000 1200.140000 365.000000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.630000 0.000000 1184.770000 0.490000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.0855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.1649 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.621 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 556.16 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1189.430000 0.000000 1189.570000 0.490000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.984 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.115 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.104 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.488 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 555.644 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1191.430000 0.000000 1191.570000 0.490000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.984 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 48.115 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.104 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.6842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 102.488 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 555.644 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1187.030000 0.000000 1187.170000 0.490000 ;
    END
  END user_irq[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 7.840000 7.680000 1192.300000 9.280000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1190.700000 7.680000 1192.300000 922.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.840000 920.960000 1192.300000 922.560000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.840000 7.680000 9.440000 922.560000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 623.410000 441.830000 625.150000 829.810000 ;
      LAYER met4 ;
        RECT 1091.930000 441.830000 1093.670000 829.810000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 109.630000 441.830000 111.370000 829.810000 ;
      LAYER met4 ;
        RECT 578.150000 441.830000 579.890000 829.810000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 4.640000 4.480000 1195.500000 6.080000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1193.900000 4.480000 1195.500000 925.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.640000 924.160000 1195.500000 925.760000 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.640000 4.480000 6.240000 925.760000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1095.330000 438.430000 1097.070000 833.210000 ;
      LAYER met4 ;
        RECT 620.010000 438.430000 621.750000 833.210000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 581.550000 438.430000 583.290000 833.210000 ;
      LAYER met4 ;
        RECT 106.230000 438.430000 107.970000 833.210000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1200.140000 930.580000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1200.140000 930.580000 ;
    #LAYER met2 ;
      RECT 1191.210000 929.950000 1200.140000 930.580000 ;
      RECT 1158.010000 929.950000 1190.790000 930.580000 ;
      RECT 1124.010000 929.950000 1157.590000 930.580000 ;
      RECT 1089.910000 929.950000 1123.590000 930.580000 ;
      RECT 1055.910000 929.950000 1089.490000 930.580000 ;
      RECT 1021.810000 929.950000 1055.490000 930.580000 ;
      RECT 987.810000 929.950000 1021.390000 930.580000 ;
      RECT 953.710000 929.950000 987.390000 930.580000 ;
      RECT 919.710000 929.950000 953.290000 930.580000 ;
      RECT 885.610000 929.950000 919.290000 930.580000 ;
      RECT 851.510000 929.950000 885.190000 930.580000 ;
      RECT 817.510000 929.950000 851.090000 930.580000 ;
      RECT 783.410000 929.950000 817.090000 930.580000 ;
      RECT 749.410000 929.950000 782.990000 930.580000 ;
      RECT 715.310000 929.950000 748.990000 930.580000 ;
      RECT 681.210000 929.950000 714.890000 930.580000 ;
      RECT 647.210000 929.950000 680.790000 930.580000 ;
      RECT 613.210000 929.950000 646.790000 930.580000 ;
      RECT 579.110000 929.950000 612.790000 930.580000 ;
      RECT 545.010000 929.950000 578.690000 930.580000 ;
      RECT 511.010000 929.950000 544.590000 930.580000 ;
      RECT 476.910000 929.950000 510.590000 930.580000 ;
      RECT 442.910000 929.950000 476.490000 930.580000 ;
      RECT 408.810000 929.950000 442.490000 930.580000 ;
      RECT 374.710000 929.950000 408.390000 930.580000 ;
      RECT 340.710000 929.950000 374.290000 930.580000 ;
      RECT 306.710000 929.950000 340.290000 930.580000 ;
      RECT 272.610000 929.950000 306.290000 930.580000 ;
      RECT 238.510000 929.950000 272.190000 930.580000 ;
      RECT 204.510000 929.950000 238.090000 930.580000 ;
      RECT 170.410000 929.950000 204.090000 930.580000 ;
      RECT 136.310000 929.950000 169.990000 930.580000 ;
      RECT 102.310000 929.950000 135.890000 930.580000 ;
      RECT 68.210000 929.950000 101.890000 930.580000 ;
      RECT 34.210000 929.950000 67.790000 930.580000 ;
      RECT 1.310000 929.950000 33.790000 930.580000 ;
      RECT 0.000000 929.950000 0.890000 930.580000 ;
      RECT 0.000000 0.630000 1200.140000 929.950000 ;
      RECT 1191.710000 0.000000 1200.140000 0.630000 ;
      RECT 1189.710000 0.000000 1191.290000 0.630000 ;
      RECT 1187.310000 0.000000 1189.290000 0.630000 ;
      RECT 1184.910000 0.000000 1186.890000 0.630000 ;
      RECT 1182.510000 0.000000 1184.490000 0.630000 ;
      RECT 1180.010000 0.000000 1182.090000 0.630000 ;
      RECT 1177.610000 0.000000 1179.590000 0.630000 ;
      RECT 1175.210000 0.000000 1177.190000 0.630000 ;
      RECT 1172.810000 0.000000 1174.790000 0.630000 ;
      RECT 1170.410000 0.000000 1172.390000 0.630000 ;
      RECT 1167.910000 0.000000 1169.990000 0.630000 ;
      RECT 1165.510000 0.000000 1167.490000 0.630000 ;
      RECT 1163.110000 0.000000 1165.090000 0.630000 ;
      RECT 1160.710000 0.000000 1162.690000 0.630000 ;
      RECT 1158.310000 0.000000 1160.290000 0.630000 ;
      RECT 1155.810000 0.000000 1157.890000 0.630000 ;
      RECT 1153.410000 0.000000 1155.390000 0.630000 ;
      RECT 1151.010000 0.000000 1152.990000 0.630000 ;
      RECT 1148.610000 0.000000 1150.590000 0.630000 ;
      RECT 1146.210000 0.000000 1148.190000 0.630000 ;
      RECT 1143.710000 0.000000 1145.790000 0.630000 ;
      RECT 1141.310000 0.000000 1143.290000 0.630000 ;
      RECT 1138.910000 0.000000 1140.890000 0.630000 ;
      RECT 1136.510000 0.000000 1138.490000 0.630000 ;
      RECT 1134.110000 0.000000 1136.090000 0.630000 ;
      RECT 1131.710000 0.000000 1133.690000 0.630000 ;
      RECT 1129.210000 0.000000 1131.290000 0.630000 ;
      RECT 1126.810000 0.000000 1128.790000 0.630000 ;
      RECT 1124.410000 0.000000 1126.390000 0.630000 ;
      RECT 1122.010000 0.000000 1123.990000 0.630000 ;
      RECT 1119.610000 0.000000 1121.590000 0.630000 ;
      RECT 1117.110000 0.000000 1119.190000 0.630000 ;
      RECT 1114.710000 0.000000 1116.690000 0.630000 ;
      RECT 1112.310000 0.000000 1114.290000 0.630000 ;
      RECT 1109.910000 0.000000 1111.890000 0.630000 ;
      RECT 1107.510000 0.000000 1109.490000 0.630000 ;
      RECT 1105.010000 0.000000 1107.090000 0.630000 ;
      RECT 1102.610000 0.000000 1104.590000 0.630000 ;
      RECT 1100.210000 0.000000 1102.190000 0.630000 ;
      RECT 1097.810000 0.000000 1099.790000 0.630000 ;
      RECT 1095.410000 0.000000 1097.390000 0.630000 ;
      RECT 1093.010000 0.000000 1094.990000 0.630000 ;
      RECT 1090.610000 0.000000 1092.590000 0.630000 ;
      RECT 1088.210000 0.000000 1090.190000 0.630000 ;
      RECT 1085.810000 0.000000 1087.790000 0.630000 ;
      RECT 1083.310000 0.000000 1085.390000 0.630000 ;
      RECT 1080.910000 0.000000 1082.890000 0.630000 ;
      RECT 1078.510000 0.000000 1080.490000 0.630000 ;
      RECT 1076.110000 0.000000 1078.090000 0.630000 ;
      RECT 1073.710000 0.000000 1075.690000 0.630000 ;
      RECT 1071.210000 0.000000 1073.290000 0.630000 ;
      RECT 1068.810000 0.000000 1070.790000 0.630000 ;
      RECT 1066.410000 0.000000 1068.390000 0.630000 ;
      RECT 1064.010000 0.000000 1065.990000 0.630000 ;
      RECT 1061.610000 0.000000 1063.590000 0.630000 ;
      RECT 1059.110000 0.000000 1061.190000 0.630000 ;
      RECT 1056.710000 0.000000 1058.690000 0.630000 ;
      RECT 1054.310000 0.000000 1056.290000 0.630000 ;
      RECT 1051.910000 0.000000 1053.890000 0.630000 ;
      RECT 1049.510000 0.000000 1051.490000 0.630000 ;
      RECT 1047.010000 0.000000 1049.090000 0.630000 ;
      RECT 1044.610000 0.000000 1046.590000 0.630000 ;
      RECT 1042.210000 0.000000 1044.190000 0.630000 ;
      RECT 1039.810000 0.000000 1041.790000 0.630000 ;
      RECT 1037.410000 0.000000 1039.390000 0.630000 ;
      RECT 1035.010000 0.000000 1036.990000 0.630000 ;
      RECT 1032.510000 0.000000 1034.590000 0.630000 ;
      RECT 1030.110000 0.000000 1032.090000 0.630000 ;
      RECT 1027.710000 0.000000 1029.690000 0.630000 ;
      RECT 1025.310000 0.000000 1027.290000 0.630000 ;
      RECT 1022.910000 0.000000 1024.890000 0.630000 ;
      RECT 1020.410000 0.000000 1022.490000 0.630000 ;
      RECT 1018.010000 0.000000 1019.990000 0.630000 ;
      RECT 1015.610000 0.000000 1017.590000 0.630000 ;
      RECT 1013.210000 0.000000 1015.190000 0.630000 ;
      RECT 1010.810000 0.000000 1012.790000 0.630000 ;
      RECT 1008.310000 0.000000 1010.390000 0.630000 ;
      RECT 1005.910000 0.000000 1007.890000 0.630000 ;
      RECT 1003.510000 0.000000 1005.490000 0.630000 ;
      RECT 1001.110000 0.000000 1003.090000 0.630000 ;
      RECT 998.710000 0.000000 1000.690000 0.630000 ;
      RECT 996.210000 0.000000 998.290000 0.630000 ;
      RECT 993.810000 0.000000 995.790000 0.630000 ;
      RECT 991.410000 0.000000 993.390000 0.630000 ;
      RECT 989.010000 0.000000 990.990000 0.630000 ;
      RECT 986.610000 0.000000 988.590000 0.630000 ;
      RECT 984.210000 0.000000 986.190000 0.630000 ;
      RECT 981.710000 0.000000 983.790000 0.630000 ;
      RECT 979.310000 0.000000 981.290000 0.630000 ;
      RECT 976.910000 0.000000 978.890000 0.630000 ;
      RECT 974.510000 0.000000 976.490000 0.630000 ;
      RECT 972.110000 0.000000 974.090000 0.630000 ;
      RECT 969.710000 0.000000 971.690000 0.630000 ;
      RECT 967.310000 0.000000 969.290000 0.630000 ;
      RECT 964.910000 0.000000 966.890000 0.630000 ;
      RECT 962.410000 0.000000 964.490000 0.630000 ;
      RECT 960.010000 0.000000 961.990000 0.630000 ;
      RECT 957.610000 0.000000 959.590000 0.630000 ;
      RECT 955.210000 0.000000 957.190000 0.630000 ;
      RECT 952.810000 0.000000 954.790000 0.630000 ;
      RECT 950.310000 0.000000 952.390000 0.630000 ;
      RECT 947.910000 0.000000 949.890000 0.630000 ;
      RECT 945.510000 0.000000 947.490000 0.630000 ;
      RECT 943.110000 0.000000 945.090000 0.630000 ;
      RECT 940.710000 0.000000 942.690000 0.630000 ;
      RECT 938.310000 0.000000 940.290000 0.630000 ;
      RECT 935.810000 0.000000 937.890000 0.630000 ;
      RECT 933.410000 0.000000 935.390000 0.630000 ;
      RECT 931.010000 0.000000 932.990000 0.630000 ;
      RECT 928.610000 0.000000 930.590000 0.630000 ;
      RECT 926.210000 0.000000 928.190000 0.630000 ;
      RECT 923.710000 0.000000 925.790000 0.630000 ;
      RECT 921.310000 0.000000 923.290000 0.630000 ;
      RECT 918.910000 0.000000 920.890000 0.630000 ;
      RECT 916.510000 0.000000 918.490000 0.630000 ;
      RECT 914.110000 0.000000 916.090000 0.630000 ;
      RECT 911.610000 0.000000 913.690000 0.630000 ;
      RECT 909.210000 0.000000 911.190000 0.630000 ;
      RECT 906.810000 0.000000 908.790000 0.630000 ;
      RECT 904.410000 0.000000 906.390000 0.630000 ;
      RECT 902.010000 0.000000 903.990000 0.630000 ;
      RECT 899.510000 0.000000 901.590000 0.630000 ;
      RECT 897.110000 0.000000 899.090000 0.630000 ;
      RECT 894.710000 0.000000 896.690000 0.630000 ;
      RECT 892.310000 0.000000 894.290000 0.630000 ;
      RECT 889.910000 0.000000 891.890000 0.630000 ;
      RECT 887.510000 0.000000 889.490000 0.630000 ;
      RECT 885.010000 0.000000 887.090000 0.630000 ;
      RECT 882.610000 0.000000 884.590000 0.630000 ;
      RECT 880.210000 0.000000 882.190000 0.630000 ;
      RECT 877.810000 0.000000 879.790000 0.630000 ;
      RECT 875.410000 0.000000 877.390000 0.630000 ;
      RECT 872.910000 0.000000 874.990000 0.630000 ;
      RECT 870.510000 0.000000 872.490000 0.630000 ;
      RECT 868.110000 0.000000 870.090000 0.630000 ;
      RECT 865.710000 0.000000 867.690000 0.630000 ;
      RECT 863.310000 0.000000 865.290000 0.630000 ;
      RECT 860.810000 0.000000 862.890000 0.630000 ;
      RECT 858.410000 0.000000 860.390000 0.630000 ;
      RECT 856.010000 0.000000 857.990000 0.630000 ;
      RECT 853.610000 0.000000 855.590000 0.630000 ;
      RECT 851.210000 0.000000 853.190000 0.630000 ;
      RECT 848.810000 0.000000 850.790000 0.630000 ;
      RECT 846.410000 0.000000 848.390000 0.630000 ;
      RECT 844.010000 0.000000 845.990000 0.630000 ;
      RECT 841.610000 0.000000 843.590000 0.630000 ;
      RECT 839.110000 0.000000 841.190000 0.630000 ;
      RECT 836.710000 0.000000 838.690000 0.630000 ;
      RECT 834.310000 0.000000 836.290000 0.630000 ;
      RECT 831.910000 0.000000 833.890000 0.630000 ;
      RECT 829.510000 0.000000 831.490000 0.630000 ;
      RECT 827.010000 0.000000 829.090000 0.630000 ;
      RECT 824.610000 0.000000 826.590000 0.630000 ;
      RECT 822.210000 0.000000 824.190000 0.630000 ;
      RECT 819.810000 0.000000 821.790000 0.630000 ;
      RECT 817.410000 0.000000 819.390000 0.630000 ;
      RECT 814.910000 0.000000 816.990000 0.630000 ;
      RECT 812.510000 0.000000 814.490000 0.630000 ;
      RECT 810.110000 0.000000 812.090000 0.630000 ;
      RECT 807.710000 0.000000 809.690000 0.630000 ;
      RECT 805.310000 0.000000 807.290000 0.630000 ;
      RECT 802.810000 0.000000 804.890000 0.630000 ;
      RECT 800.410000 0.000000 802.390000 0.630000 ;
      RECT 798.010000 0.000000 799.990000 0.630000 ;
      RECT 795.610000 0.000000 797.590000 0.630000 ;
      RECT 793.210000 0.000000 795.190000 0.630000 ;
      RECT 790.810000 0.000000 792.790000 0.630000 ;
      RECT 788.310000 0.000000 790.390000 0.630000 ;
      RECT 785.910000 0.000000 787.890000 0.630000 ;
      RECT 783.510000 0.000000 785.490000 0.630000 ;
      RECT 781.110000 0.000000 783.090000 0.630000 ;
      RECT 778.710000 0.000000 780.690000 0.630000 ;
      RECT 776.210000 0.000000 778.290000 0.630000 ;
      RECT 773.810000 0.000000 775.790000 0.630000 ;
      RECT 771.410000 0.000000 773.390000 0.630000 ;
      RECT 769.010000 0.000000 770.990000 0.630000 ;
      RECT 766.610000 0.000000 768.590000 0.630000 ;
      RECT 764.110000 0.000000 766.190000 0.630000 ;
      RECT 761.710000 0.000000 763.690000 0.630000 ;
      RECT 759.310000 0.000000 761.290000 0.630000 ;
      RECT 756.910000 0.000000 758.890000 0.630000 ;
      RECT 754.510000 0.000000 756.490000 0.630000 ;
      RECT 752.010000 0.000000 754.090000 0.630000 ;
      RECT 749.610000 0.000000 751.590000 0.630000 ;
      RECT 747.210000 0.000000 749.190000 0.630000 ;
      RECT 744.810000 0.000000 746.790000 0.630000 ;
      RECT 742.410000 0.000000 744.390000 0.630000 ;
      RECT 740.010000 0.000000 741.990000 0.630000 ;
      RECT 737.510000 0.000000 739.590000 0.630000 ;
      RECT 735.110000 0.000000 737.090000 0.630000 ;
      RECT 732.710000 0.000000 734.690000 0.630000 ;
      RECT 730.310000 0.000000 732.290000 0.630000 ;
      RECT 727.910000 0.000000 729.890000 0.630000 ;
      RECT 725.510000 0.000000 727.490000 0.630000 ;
      RECT 723.110000 0.000000 725.090000 0.630000 ;
      RECT 720.710000 0.000000 722.690000 0.630000 ;
      RECT 718.210000 0.000000 720.290000 0.630000 ;
      RECT 715.810000 0.000000 717.790000 0.630000 ;
      RECT 713.410000 0.000000 715.390000 0.630000 ;
      RECT 711.010000 0.000000 712.990000 0.630000 ;
      RECT 708.610000 0.000000 710.590000 0.630000 ;
      RECT 706.110000 0.000000 708.190000 0.630000 ;
      RECT 703.710000 0.000000 705.690000 0.630000 ;
      RECT 701.310000 0.000000 703.290000 0.630000 ;
      RECT 698.910000 0.000000 700.890000 0.630000 ;
      RECT 696.510000 0.000000 698.490000 0.630000 ;
      RECT 694.110000 0.000000 696.090000 0.630000 ;
      RECT 691.610000 0.000000 693.690000 0.630000 ;
      RECT 689.210000 0.000000 691.190000 0.630000 ;
      RECT 686.810000 0.000000 688.790000 0.630000 ;
      RECT 684.410000 0.000000 686.390000 0.630000 ;
      RECT 682.010000 0.000000 683.990000 0.630000 ;
      RECT 679.510000 0.000000 681.590000 0.630000 ;
      RECT 677.110000 0.000000 679.090000 0.630000 ;
      RECT 674.710000 0.000000 676.690000 0.630000 ;
      RECT 672.310000 0.000000 674.290000 0.630000 ;
      RECT 669.910000 0.000000 671.890000 0.630000 ;
      RECT 667.410000 0.000000 669.490000 0.630000 ;
      RECT 665.010000 0.000000 666.990000 0.630000 ;
      RECT 662.610000 0.000000 664.590000 0.630000 ;
      RECT 660.210000 0.000000 662.190000 0.630000 ;
      RECT 657.810000 0.000000 659.790000 0.630000 ;
      RECT 655.310000 0.000000 657.390000 0.630000 ;
      RECT 652.910000 0.000000 654.890000 0.630000 ;
      RECT 650.510000 0.000000 652.490000 0.630000 ;
      RECT 648.110000 0.000000 650.090000 0.630000 ;
      RECT 645.710000 0.000000 647.690000 0.630000 ;
      RECT 643.310000 0.000000 645.290000 0.630000 ;
      RECT 640.810000 0.000000 642.890000 0.630000 ;
      RECT 638.410000 0.000000 640.390000 0.630000 ;
      RECT 636.010000 0.000000 637.990000 0.630000 ;
      RECT 633.610000 0.000000 635.590000 0.630000 ;
      RECT 631.210000 0.000000 633.190000 0.630000 ;
      RECT 628.710000 0.000000 630.790000 0.630000 ;
      RECT 626.310000 0.000000 628.290000 0.630000 ;
      RECT 623.910000 0.000000 625.890000 0.630000 ;
      RECT 621.510000 0.000000 623.490000 0.630000 ;
      RECT 619.110000 0.000000 621.090000 0.630000 ;
      RECT 616.610000 0.000000 618.690000 0.630000 ;
      RECT 614.210000 0.000000 616.190000 0.630000 ;
      RECT 611.810000 0.000000 613.790000 0.630000 ;
      RECT 609.410000 0.000000 611.390000 0.630000 ;
      RECT 607.010000 0.000000 608.990000 0.630000 ;
      RECT 604.610000 0.000000 606.590000 0.630000 ;
      RECT 602.210000 0.000000 604.190000 0.630000 ;
      RECT 599.810000 0.000000 601.790000 0.630000 ;
      RECT 597.410000 0.000000 599.390000 0.630000 ;
      RECT 594.910000 0.000000 596.990000 0.630000 ;
      RECT 592.510000 0.000000 594.490000 0.630000 ;
      RECT 590.110000 0.000000 592.090000 0.630000 ;
      RECT 587.710000 0.000000 589.690000 0.630000 ;
      RECT 585.310000 0.000000 587.290000 0.630000 ;
      RECT 582.810000 0.000000 584.890000 0.630000 ;
      RECT 580.410000 0.000000 582.390000 0.630000 ;
      RECT 578.010000 0.000000 579.990000 0.630000 ;
      RECT 575.610000 0.000000 577.590000 0.630000 ;
      RECT 573.210000 0.000000 575.190000 0.630000 ;
      RECT 570.710000 0.000000 572.790000 0.630000 ;
      RECT 568.310000 0.000000 570.290000 0.630000 ;
      RECT 565.910000 0.000000 567.890000 0.630000 ;
      RECT 563.510000 0.000000 565.490000 0.630000 ;
      RECT 561.110000 0.000000 563.090000 0.630000 ;
      RECT 558.610000 0.000000 560.690000 0.630000 ;
      RECT 556.210000 0.000000 558.190000 0.630000 ;
      RECT 553.810000 0.000000 555.790000 0.630000 ;
      RECT 551.410000 0.000000 553.390000 0.630000 ;
      RECT 549.010000 0.000000 550.990000 0.630000 ;
      RECT 546.610000 0.000000 548.590000 0.630000 ;
      RECT 544.110000 0.000000 546.190000 0.630000 ;
      RECT 541.710000 0.000000 543.690000 0.630000 ;
      RECT 539.310000 0.000000 541.290000 0.630000 ;
      RECT 536.910000 0.000000 538.890000 0.630000 ;
      RECT 534.510000 0.000000 536.490000 0.630000 ;
      RECT 532.010000 0.000000 534.090000 0.630000 ;
      RECT 529.610000 0.000000 531.590000 0.630000 ;
      RECT 527.210000 0.000000 529.190000 0.630000 ;
      RECT 524.810000 0.000000 526.790000 0.630000 ;
      RECT 522.410000 0.000000 524.390000 0.630000 ;
      RECT 519.910000 0.000000 521.990000 0.630000 ;
      RECT 517.510000 0.000000 519.490000 0.630000 ;
      RECT 515.110000 0.000000 517.090000 0.630000 ;
      RECT 512.710000 0.000000 514.690000 0.630000 ;
      RECT 510.310000 0.000000 512.290000 0.630000 ;
      RECT 507.810000 0.000000 509.890000 0.630000 ;
      RECT 505.410000 0.000000 507.390000 0.630000 ;
      RECT 503.010000 0.000000 504.990000 0.630000 ;
      RECT 500.610000 0.000000 502.590000 0.630000 ;
      RECT 498.210000 0.000000 500.190000 0.630000 ;
      RECT 495.810000 0.000000 497.790000 0.630000 ;
      RECT 493.310000 0.000000 495.390000 0.630000 ;
      RECT 490.910000 0.000000 492.890000 0.630000 ;
      RECT 488.510000 0.000000 490.490000 0.630000 ;
      RECT 486.110000 0.000000 488.090000 0.630000 ;
      RECT 483.710000 0.000000 485.690000 0.630000 ;
      RECT 481.310000 0.000000 483.290000 0.630000 ;
      RECT 478.910000 0.000000 480.890000 0.630000 ;
      RECT 476.510000 0.000000 478.490000 0.630000 ;
      RECT 474.010000 0.000000 476.090000 0.630000 ;
      RECT 471.610000 0.000000 473.590000 0.630000 ;
      RECT 469.210000 0.000000 471.190000 0.630000 ;
      RECT 466.810000 0.000000 468.790000 0.630000 ;
      RECT 464.410000 0.000000 466.390000 0.630000 ;
      RECT 461.910000 0.000000 463.990000 0.630000 ;
      RECT 459.510000 0.000000 461.490000 0.630000 ;
      RECT 457.110000 0.000000 459.090000 0.630000 ;
      RECT 454.710000 0.000000 456.690000 0.630000 ;
      RECT 452.310000 0.000000 454.290000 0.630000 ;
      RECT 449.910000 0.000000 451.890000 0.630000 ;
      RECT 447.410000 0.000000 449.490000 0.630000 ;
      RECT 445.010000 0.000000 446.990000 0.630000 ;
      RECT 442.610000 0.000000 444.590000 0.630000 ;
      RECT 440.210000 0.000000 442.190000 0.630000 ;
      RECT 437.810000 0.000000 439.790000 0.630000 ;
      RECT 435.310000 0.000000 437.390000 0.630000 ;
      RECT 432.910000 0.000000 434.890000 0.630000 ;
      RECT 430.510000 0.000000 432.490000 0.630000 ;
      RECT 428.110000 0.000000 430.090000 0.630000 ;
      RECT 425.710000 0.000000 427.690000 0.630000 ;
      RECT 423.210000 0.000000 425.290000 0.630000 ;
      RECT 420.810000 0.000000 422.790000 0.630000 ;
      RECT 418.410000 0.000000 420.390000 0.630000 ;
      RECT 416.010000 0.000000 417.990000 0.630000 ;
      RECT 413.610000 0.000000 415.590000 0.630000 ;
      RECT 411.110000 0.000000 413.190000 0.630000 ;
      RECT 408.710000 0.000000 410.690000 0.630000 ;
      RECT 406.310000 0.000000 408.290000 0.630000 ;
      RECT 403.910000 0.000000 405.890000 0.630000 ;
      RECT 401.510000 0.000000 403.490000 0.630000 ;
      RECT 399.110000 0.000000 401.090000 0.630000 ;
      RECT 396.610000 0.000000 398.690000 0.630000 ;
      RECT 394.210000 0.000000 396.190000 0.630000 ;
      RECT 391.810000 0.000000 393.790000 0.630000 ;
      RECT 389.410000 0.000000 391.390000 0.630000 ;
      RECT 387.010000 0.000000 388.990000 0.630000 ;
      RECT 384.510000 0.000000 386.590000 0.630000 ;
      RECT 382.110000 0.000000 384.090000 0.630000 ;
      RECT 379.710000 0.000000 381.690000 0.630000 ;
      RECT 377.310000 0.000000 379.290000 0.630000 ;
      RECT 374.910000 0.000000 376.890000 0.630000 ;
      RECT 372.410000 0.000000 374.490000 0.630000 ;
      RECT 370.010000 0.000000 371.990000 0.630000 ;
      RECT 367.610000 0.000000 369.590000 0.630000 ;
      RECT 365.210000 0.000000 367.190000 0.630000 ;
      RECT 362.810000 0.000000 364.790000 0.630000 ;
      RECT 360.410000 0.000000 362.390000 0.630000 ;
      RECT 358.010000 0.000000 359.990000 0.630000 ;
      RECT 355.610000 0.000000 357.590000 0.630000 ;
      RECT 353.110000 0.000000 355.190000 0.630000 ;
      RECT 350.710000 0.000000 352.690000 0.630000 ;
      RECT 348.310000 0.000000 350.290000 0.630000 ;
      RECT 345.910000 0.000000 347.890000 0.630000 ;
      RECT 343.510000 0.000000 345.490000 0.630000 ;
      RECT 341.110000 0.000000 343.090000 0.630000 ;
      RECT 338.610000 0.000000 340.690000 0.630000 ;
      RECT 336.210000 0.000000 338.190000 0.630000 ;
      RECT 333.810000 0.000000 335.790000 0.630000 ;
      RECT 331.410000 0.000000 333.390000 0.630000 ;
      RECT 329.010000 0.000000 330.990000 0.630000 ;
      RECT 326.510000 0.000000 328.590000 0.630000 ;
      RECT 324.110000 0.000000 326.090000 0.630000 ;
      RECT 321.710000 0.000000 323.690000 0.630000 ;
      RECT 319.310000 0.000000 321.290000 0.630000 ;
      RECT 316.910000 0.000000 318.890000 0.630000 ;
      RECT 314.410000 0.000000 316.490000 0.630000 ;
      RECT 312.010000 0.000000 313.990000 0.630000 ;
      RECT 309.610000 0.000000 311.590000 0.630000 ;
      RECT 307.210000 0.000000 309.190000 0.630000 ;
      RECT 304.810000 0.000000 306.790000 0.630000 ;
      RECT 302.410000 0.000000 304.390000 0.630000 ;
      RECT 299.910000 0.000000 301.990000 0.630000 ;
      RECT 297.510000 0.000000 299.490000 0.630000 ;
      RECT 295.110000 0.000000 297.090000 0.630000 ;
      RECT 292.710000 0.000000 294.690000 0.630000 ;
      RECT 290.310000 0.000000 292.290000 0.630000 ;
      RECT 287.810000 0.000000 289.890000 0.630000 ;
      RECT 285.410000 0.000000 287.390000 0.630000 ;
      RECT 283.010000 0.000000 284.990000 0.630000 ;
      RECT 280.610000 0.000000 282.590000 0.630000 ;
      RECT 278.210000 0.000000 280.190000 0.630000 ;
      RECT 275.710000 0.000000 277.790000 0.630000 ;
      RECT 273.310000 0.000000 275.290000 0.630000 ;
      RECT 270.910000 0.000000 272.890000 0.630000 ;
      RECT 268.510000 0.000000 270.490000 0.630000 ;
      RECT 266.110000 0.000000 268.090000 0.630000 ;
      RECT 263.610000 0.000000 265.690000 0.630000 ;
      RECT 261.210000 0.000000 263.190000 0.630000 ;
      RECT 258.810000 0.000000 260.790000 0.630000 ;
      RECT 256.410000 0.000000 258.390000 0.630000 ;
      RECT 254.010000 0.000000 255.990000 0.630000 ;
      RECT 251.610000 0.000000 253.590000 0.630000 ;
      RECT 249.110000 0.000000 251.190000 0.630000 ;
      RECT 246.710000 0.000000 248.690000 0.630000 ;
      RECT 244.410000 0.000000 246.290000 0.630000 ;
      RECT 241.910000 0.000000 243.990000 0.630000 ;
      RECT 239.510000 0.000000 241.490000 0.630000 ;
      RECT 237.110000 0.000000 239.090000 0.630000 ;
      RECT 234.710000 0.000000 236.690000 0.630000 ;
      RECT 232.310000 0.000000 234.290000 0.630000 ;
      RECT 229.810000 0.000000 231.890000 0.630000 ;
      RECT 227.410000 0.000000 229.390000 0.630000 ;
      RECT 225.010000 0.000000 226.990000 0.630000 ;
      RECT 222.610000 0.000000 224.590000 0.630000 ;
      RECT 220.210000 0.000000 222.190000 0.630000 ;
      RECT 217.710000 0.000000 219.790000 0.630000 ;
      RECT 215.310000 0.000000 217.290000 0.630000 ;
      RECT 212.910000 0.000000 214.890000 0.630000 ;
      RECT 210.510000 0.000000 212.490000 0.630000 ;
      RECT 208.110000 0.000000 210.090000 0.630000 ;
      RECT 205.610000 0.000000 207.690000 0.630000 ;
      RECT 203.210000 0.000000 205.190000 0.630000 ;
      RECT 200.810000 0.000000 202.790000 0.630000 ;
      RECT 198.410000 0.000000 200.390000 0.630000 ;
      RECT 196.010000 0.000000 197.990000 0.630000 ;
      RECT 193.610000 0.000000 195.590000 0.630000 ;
      RECT 191.110000 0.000000 193.190000 0.630000 ;
      RECT 188.710000 0.000000 190.690000 0.630000 ;
      RECT 186.310000 0.000000 188.290000 0.630000 ;
      RECT 183.910000 0.000000 185.890000 0.630000 ;
      RECT 181.510000 0.000000 183.490000 0.630000 ;
      RECT 179.010000 0.000000 181.090000 0.630000 ;
      RECT 176.610000 0.000000 178.590000 0.630000 ;
      RECT 174.210000 0.000000 176.190000 0.630000 ;
      RECT 171.810000 0.000000 173.790000 0.630000 ;
      RECT 169.410000 0.000000 171.390000 0.630000 ;
      RECT 166.910000 0.000000 168.990000 0.630000 ;
      RECT 164.510000 0.000000 166.490000 0.630000 ;
      RECT 162.110000 0.000000 164.090000 0.630000 ;
      RECT 159.710000 0.000000 161.690000 0.630000 ;
      RECT 157.310000 0.000000 159.290000 0.630000 ;
      RECT 154.910000 0.000000 156.890000 0.630000 ;
      RECT 152.410000 0.000000 154.490000 0.630000 ;
      RECT 150.010000 0.000000 151.990000 0.630000 ;
      RECT 147.610000 0.000000 149.590000 0.630000 ;
      RECT 145.210000 0.000000 147.190000 0.630000 ;
      RECT 142.810000 0.000000 144.790000 0.630000 ;
      RECT 140.310000 0.000000 142.390000 0.630000 ;
      RECT 137.910000 0.000000 139.890000 0.630000 ;
      RECT 135.510000 0.000000 137.490000 0.630000 ;
      RECT 133.110000 0.000000 135.090000 0.630000 ;
      RECT 130.710000 0.000000 132.690000 0.630000 ;
      RECT 128.210000 0.000000 130.290000 0.630000 ;
      RECT 125.810000 0.000000 127.790000 0.630000 ;
      RECT 123.510000 0.000000 125.390000 0.630000 ;
      RECT 121.010000 0.000000 123.090000 0.630000 ;
      RECT 118.610000 0.000000 120.590000 0.630000 ;
      RECT 116.210000 0.000000 118.190000 0.630000 ;
      RECT 113.810000 0.000000 115.790000 0.630000 ;
      RECT 111.410000 0.000000 113.390000 0.630000 ;
      RECT 108.910000 0.000000 110.990000 0.630000 ;
      RECT 106.510000 0.000000 108.490000 0.630000 ;
      RECT 104.110000 0.000000 106.090000 0.630000 ;
      RECT 101.710000 0.000000 103.690000 0.630000 ;
      RECT 99.310000 0.000000 101.290000 0.630000 ;
      RECT 96.910000 0.000000 98.890000 0.630000 ;
      RECT 94.410000 0.000000 96.490000 0.630000 ;
      RECT 92.010000 0.000000 93.990000 0.630000 ;
      RECT 89.610000 0.000000 91.590000 0.630000 ;
      RECT 87.210000 0.000000 89.190000 0.630000 ;
      RECT 84.810000 0.000000 86.790000 0.630000 ;
      RECT 82.310000 0.000000 84.390000 0.630000 ;
      RECT 79.910000 0.000000 81.890000 0.630000 ;
      RECT 77.510000 0.000000 79.490000 0.630000 ;
      RECT 75.110000 0.000000 77.090000 0.630000 ;
      RECT 72.710000 0.000000 74.690000 0.630000 ;
      RECT 70.210000 0.000000 72.290000 0.630000 ;
      RECT 67.810000 0.000000 69.790000 0.630000 ;
      RECT 65.410000 0.000000 67.390000 0.630000 ;
      RECT 63.010000 0.000000 64.990000 0.630000 ;
      RECT 60.610000 0.000000 62.590000 0.630000 ;
      RECT 58.110000 0.000000 60.190000 0.630000 ;
      RECT 55.710000 0.000000 57.690000 0.630000 ;
      RECT 53.310000 0.000000 55.290000 0.630000 ;
      RECT 50.910000 0.000000 52.890000 0.630000 ;
      RECT 48.510000 0.000000 50.490000 0.630000 ;
      RECT 46.110000 0.000000 48.090000 0.630000 ;
      RECT 43.610000 0.000000 45.690000 0.630000 ;
      RECT 41.210000 0.000000 43.190000 0.630000 ;
      RECT 38.810000 0.000000 40.790000 0.630000 ;
      RECT 36.410000 0.000000 38.390000 0.630000 ;
      RECT 34.010000 0.000000 35.990000 0.630000 ;
      RECT 31.510000 0.000000 33.590000 0.630000 ;
      RECT 29.110000 0.000000 31.090000 0.630000 ;
      RECT 26.710000 0.000000 28.690000 0.630000 ;
      RECT 24.310000 0.000000 26.290000 0.630000 ;
      RECT 21.910000 0.000000 23.890000 0.630000 ;
      RECT 19.410000 0.000000 21.490000 0.630000 ;
      RECT 17.010000 0.000000 18.990000 0.630000 ;
      RECT 14.610000 0.000000 16.590000 0.630000 ;
      RECT 12.210000 0.000000 14.190000 0.630000 ;
      RECT 9.810000 0.000000 11.790000 0.630000 ;
      RECT 7.410000 0.000000 9.390000 0.630000 ;
      RECT 4.910000 0.000000 6.990000 0.630000 ;
      RECT 2.610000 0.000000 4.490000 0.630000 ;
      RECT 0.000000 0.000000 2.190000 0.630000 ;
   # LAYER met3 ;
      RECT 0.000000 926.060000 1200.140000 930.580000 ;
      RECT 1195.800000 923.860000 1200.140000 926.060000 ;
      RECT 0.000000 923.860000 4.340000 926.060000 ;
      RECT 0.000000 922.860000 1200.140000 923.860000 ;
      RECT 1192.600000 920.660000 1200.140000 922.860000 ;
      RECT 0.000000 920.660000 7.540000 922.860000 ;
      RECT 0.000000 905.150000 1200.140000 920.660000 ;
      RECT 1.100000 904.540000 1200.140000 905.150000 ;
      RECT 1.100000 904.250000 1199.040000 904.540000 ;
      RECT 0.000000 903.640000 1199.040000 904.250000 ;
      RECT 0.000000 888.070000 1200.140000 903.640000 ;
      RECT 1.100000 887.460000 1200.140000 888.070000 ;
      RECT 1.100000 887.170000 1199.040000 887.460000 ;
      RECT 0.000000 886.560000 1199.040000 887.170000 ;
      RECT 0.000000 871.600000 1200.140000 886.560000 ;
      RECT 1.100000 870.700000 1200.140000 871.600000 ;
      RECT 0.000000 869.770000 1200.140000 870.700000 ;
      RECT 0.000000 868.870000 1199.040000 869.770000 ;
      RECT 0.000000 854.520000 1200.140000 868.870000 ;
      RECT 1.100000 853.620000 1200.140000 854.520000 ;
      RECT 0.000000 852.690000 1200.140000 853.620000 ;
      RECT 0.000000 851.790000 1199.040000 852.690000 ;
      RECT 0.000000 837.440000 1200.140000 851.790000 ;
      RECT 1.100000 836.540000 1200.140000 837.440000 ;
      RECT 0.000000 835.000000 1200.140000 836.540000 ;
      RECT 0.000000 834.100000 1199.040000 835.000000 ;
      RECT 0.000000 820.360000 1200.140000 834.100000 ;
      RECT 1.100000 819.460000 1200.140000 820.360000 ;
      RECT 0.000000 817.920000 1200.140000 819.460000 ;
      RECT 0.000000 817.020000 1199.040000 817.920000 ;
      RECT 0.000000 802.670000 1200.140000 817.020000 ;
      RECT 1.100000 801.770000 1200.140000 802.670000 ;
      RECT 0.000000 800.230000 1200.140000 801.770000 ;
      RECT 0.000000 799.330000 1199.040000 800.230000 ;
      RECT 0.000000 786.200000 1200.140000 799.330000 ;
      RECT 1.100000 785.300000 1200.140000 786.200000 ;
      RECT 0.000000 783.150000 1200.140000 785.300000 ;
      RECT 0.000000 782.250000 1199.040000 783.150000 ;
      RECT 0.000000 769.120000 1200.140000 782.250000 ;
      RECT 1.100000 768.220000 1200.140000 769.120000 ;
      RECT 0.000000 765.460000 1200.140000 768.220000 ;
      RECT 0.000000 764.560000 1199.040000 765.460000 ;
      RECT 0.000000 752.040000 1200.140000 764.560000 ;
      RECT 1.100000 751.140000 1200.140000 752.040000 ;
      RECT 0.000000 748.380000 1200.140000 751.140000 ;
      RECT 0.000000 747.480000 1199.040000 748.380000 ;
      RECT 0.000000 734.960000 1200.140000 747.480000 ;
      RECT 1.100000 734.060000 1200.140000 734.960000 ;
      RECT 0.000000 730.690000 1200.140000 734.060000 ;
      RECT 0.000000 729.790000 1199.040000 730.690000 ;
      RECT 0.000000 717.880000 1200.140000 729.790000 ;
      RECT 1.100000 716.980000 1200.140000 717.880000 ;
      RECT 0.000000 713.610000 1200.140000 716.980000 ;
      RECT 0.000000 712.710000 1199.040000 713.610000 ;
      RECT 0.000000 700.800000 1200.140000 712.710000 ;
      RECT 1.100000 699.900000 1200.140000 700.800000 ;
      RECT 0.000000 695.920000 1200.140000 699.900000 ;
      RECT 0.000000 695.020000 1199.040000 695.920000 ;
      RECT 0.000000 683.720000 1200.140000 695.020000 ;
      RECT 1.100000 682.820000 1200.140000 683.720000 ;
      RECT 0.000000 678.840000 1200.140000 682.820000 ;
      RECT 0.000000 677.940000 1199.040000 678.840000 ;
      RECT 0.000000 666.640000 1200.140000 677.940000 ;
      RECT 1.100000 665.740000 1200.140000 666.640000 ;
      RECT 0.000000 661.150000 1200.140000 665.740000 ;
      RECT 0.000000 660.250000 1199.040000 661.150000 ;
      RECT 0.000000 649.560000 1200.140000 660.250000 ;
      RECT 1.100000 648.660000 1200.140000 649.560000 ;
      RECT 0.000000 644.070000 1200.140000 648.660000 ;
      RECT 0.000000 643.170000 1199.040000 644.070000 ;
      RECT 0.000000 632.480000 1200.140000 643.170000 ;
      RECT 1.100000 631.580000 1200.140000 632.480000 ;
      RECT 0.000000 626.380000 1200.140000 631.580000 ;
      RECT 0.000000 625.480000 1199.040000 626.380000 ;
      RECT 0.000000 615.400000 1200.140000 625.480000 ;
      RECT 1.100000 614.500000 1200.140000 615.400000 ;
      RECT 0.000000 609.300000 1200.140000 614.500000 ;
      RECT 0.000000 608.400000 1199.040000 609.300000 ;
      RECT 0.000000 598.320000 1200.140000 608.400000 ;
      RECT 1.100000 597.420000 1200.140000 598.320000 ;
      RECT 0.000000 591.610000 1200.140000 597.420000 ;
      RECT 0.000000 590.710000 1199.040000 591.610000 ;
      RECT 0.000000 581.240000 1200.140000 590.710000 ;
      RECT 1.100000 580.340000 1200.140000 581.240000 ;
      RECT 0.000000 574.530000 1200.140000 580.340000 ;
      RECT 0.000000 573.630000 1199.040000 574.530000 ;
      RECT 0.000000 564.160000 1200.140000 573.630000 ;
      RECT 1.100000 563.260000 1200.140000 564.160000 ;
      RECT 0.000000 556.840000 1200.140000 563.260000 ;
      RECT 0.000000 555.940000 1199.040000 556.840000 ;
      RECT 0.000000 547.080000 1200.140000 555.940000 ;
      RECT 1.100000 546.180000 1200.140000 547.080000 ;
      RECT 0.000000 539.150000 1200.140000 546.180000 ;
      RECT 0.000000 538.250000 1199.040000 539.150000 ;
      RECT 0.000000 530.000000 1200.140000 538.250000 ;
      RECT 1.100000 529.100000 1200.140000 530.000000 ;
      RECT 0.000000 522.070000 1200.140000 529.100000 ;
      RECT 0.000000 521.170000 1199.040000 522.070000 ;
      RECT 0.000000 512.920000 1200.140000 521.170000 ;
      RECT 1.100000 512.020000 1200.140000 512.920000 ;
      RECT 0.000000 504.380000 1200.140000 512.020000 ;
      RECT 0.000000 503.480000 1199.040000 504.380000 ;
      RECT 0.000000 495.840000 1200.140000 503.480000 ;
      RECT 1.100000 494.940000 1200.140000 495.840000 ;
      RECT 0.000000 487.300000 1200.140000 494.940000 ;
      RECT 0.000000 486.400000 1199.040000 487.300000 ;
      RECT 0.000000 478.760000 1200.140000 486.400000 ;
      RECT 1.100000 477.860000 1200.140000 478.760000 ;
      RECT 0.000000 469.610000 1200.140000 477.860000 ;
      RECT 0.000000 468.710000 1199.040000 469.610000 ;
      RECT 0.000000 461.680000 1200.140000 468.710000 ;
      RECT 1.100000 460.780000 1200.140000 461.680000 ;
      RECT 0.000000 452.530000 1200.140000 460.780000 ;
      RECT 0.000000 451.630000 1199.040000 452.530000 ;
      RECT 0.000000 444.600000 1200.140000 451.630000 ;
      RECT 1.100000 443.700000 1200.140000 444.600000 ;
      RECT 0.000000 434.840000 1200.140000 443.700000 ;
      RECT 0.000000 433.940000 1199.040000 434.840000 ;
      RECT 0.000000 427.520000 1200.140000 433.940000 ;
      RECT 1.100000 426.620000 1200.140000 427.520000 ;
      RECT 0.000000 417.760000 1200.140000 426.620000 ;
      RECT 0.000000 416.860000 1199.040000 417.760000 ;
      RECT 0.000000 410.440000 1200.140000 416.860000 ;
      RECT 1.100000 409.540000 1200.140000 410.440000 ;
      RECT 0.000000 400.070000 1200.140000 409.540000 ;
      RECT 0.000000 399.170000 1199.040000 400.070000 ;
      RECT 0.000000 393.360000 1200.140000 399.170000 ;
      RECT 1.100000 392.460000 1200.140000 393.360000 ;
      RECT 0.000000 382.990000 1200.140000 392.460000 ;
      RECT 0.000000 382.090000 1199.040000 382.990000 ;
      RECT 0.000000 376.280000 1200.140000 382.090000 ;
      RECT 1.100000 375.380000 1200.140000 376.280000 ;
      RECT 0.000000 365.300000 1200.140000 375.380000 ;
      RECT 0.000000 364.400000 1199.040000 365.300000 ;
      RECT 0.000000 359.200000 1200.140000 364.400000 ;
      RECT 1.100000 358.300000 1200.140000 359.200000 ;
      RECT 0.000000 348.220000 1200.140000 358.300000 ;
      RECT 0.000000 347.320000 1199.040000 348.220000 ;
      RECT 0.000000 342.120000 1200.140000 347.320000 ;
      RECT 1.100000 341.220000 1200.140000 342.120000 ;
      RECT 0.000000 330.530000 1200.140000 341.220000 ;
      RECT 0.000000 329.630000 1199.040000 330.530000 ;
      RECT 0.000000 325.040000 1200.140000 329.630000 ;
      RECT 1.100000 324.140000 1200.140000 325.040000 ;
      RECT 0.000000 313.450000 1200.140000 324.140000 ;
      RECT 0.000000 312.550000 1199.040000 313.450000 ;
      RECT 0.000000 307.960000 1200.140000 312.550000 ;
      RECT 1.100000 307.060000 1200.140000 307.960000 ;
      RECT 0.000000 295.760000 1200.140000 307.060000 ;
      RECT 0.000000 294.860000 1199.040000 295.760000 ;
      RECT 0.000000 290.880000 1200.140000 294.860000 ;
      RECT 1.100000 289.980000 1200.140000 290.880000 ;
      RECT 0.000000 278.680000 1200.140000 289.980000 ;
      RECT 0.000000 277.780000 1199.040000 278.680000 ;
      RECT 0.000000 273.800000 1200.140000 277.780000 ;
      RECT 1.100000 272.900000 1200.140000 273.800000 ;
      RECT 0.000000 260.990000 1200.140000 272.900000 ;
      RECT 0.000000 260.090000 1199.040000 260.990000 ;
      RECT 0.000000 256.720000 1200.140000 260.090000 ;
      RECT 1.100000 255.820000 1200.140000 256.720000 ;
      RECT 0.000000 243.910000 1200.140000 255.820000 ;
      RECT 0.000000 243.010000 1199.040000 243.910000 ;
      RECT 0.000000 239.640000 1200.140000 243.010000 ;
      RECT 1.100000 238.740000 1200.140000 239.640000 ;
      RECT 0.000000 226.220000 1200.140000 238.740000 ;
      RECT 0.000000 225.320000 1199.040000 226.220000 ;
      RECT 0.000000 222.560000 1200.140000 225.320000 ;
      RECT 1.100000 221.660000 1200.140000 222.560000 ;
      RECT 0.000000 209.140000 1200.140000 221.660000 ;
      RECT 0.000000 208.240000 1199.040000 209.140000 ;
      RECT 0.000000 205.480000 1200.140000 208.240000 ;
      RECT 1.100000 204.580000 1200.140000 205.480000 ;
      RECT 0.000000 191.450000 1200.140000 204.580000 ;
      RECT 0.000000 190.550000 1199.040000 191.450000 ;
      RECT 0.000000 188.400000 1200.140000 190.550000 ;
      RECT 1.100000 187.500000 1200.140000 188.400000 ;
      RECT 0.000000 173.760000 1200.140000 187.500000 ;
      RECT 0.000000 172.860000 1199.040000 173.760000 ;
      RECT 0.000000 171.320000 1200.140000 172.860000 ;
      RECT 1.100000 170.420000 1200.140000 171.320000 ;
      RECT 0.000000 156.680000 1200.140000 170.420000 ;
      RECT 0.000000 155.780000 1199.040000 156.680000 ;
      RECT 0.000000 154.240000 1200.140000 155.780000 ;
      RECT 1.100000 153.340000 1200.140000 154.240000 ;
      RECT 0.000000 138.990000 1200.140000 153.340000 ;
      RECT 0.000000 138.090000 1199.040000 138.990000 ;
      RECT 0.000000 137.160000 1200.140000 138.090000 ;
      RECT 1.100000 136.260000 1200.140000 137.160000 ;
      RECT 0.000000 121.910000 1200.140000 136.260000 ;
      RECT 0.000000 121.010000 1199.040000 121.910000 ;
      RECT 0.000000 120.080000 1200.140000 121.010000 ;
      RECT 1.100000 119.180000 1200.140000 120.080000 ;
      RECT 0.000000 104.220000 1200.140000 119.180000 ;
      RECT 0.000000 103.320000 1199.040000 104.220000 ;
      RECT 0.000000 103.000000 1200.140000 103.320000 ;
      RECT 1.100000 102.100000 1200.140000 103.000000 ;
      RECT 0.000000 87.140000 1200.140000 102.100000 ;
      RECT 0.000000 86.240000 1199.040000 87.140000 ;
      RECT 0.000000 85.920000 1200.140000 86.240000 ;
      RECT 1.100000 85.020000 1200.140000 85.920000 ;
      RECT 0.000000 69.450000 1200.140000 85.020000 ;
      RECT 0.000000 68.840000 1199.040000 69.450000 ;
      RECT 1.100000 68.550000 1199.040000 68.840000 ;
      RECT 1.100000 67.940000 1200.140000 68.550000 ;
      RECT 0.000000 52.370000 1200.140000 67.940000 ;
      RECT 0.000000 51.760000 1199.040000 52.370000 ;
      RECT 1.100000 51.470000 1199.040000 51.760000 ;
      RECT 1.100000 50.860000 1200.140000 51.470000 ;
      RECT 0.000000 34.680000 1200.140000 50.860000 ;
      RECT 1.100000 33.780000 1199.040000 34.680000 ;
      RECT 0.000000 17.600000 1200.140000 33.780000 ;
      RECT 1.100000 16.700000 1199.040000 17.600000 ;
      RECT 0.000000 9.580000 1200.140000 16.700000 ;
      RECT 1192.600000 7.380000 1200.140000 9.580000 ;
      RECT 0.000000 7.380000 7.540000 9.580000 ;
      RECT 0.000000 6.380000 1200.140000 7.380000 ;
      RECT 1195.800000 4.180000 1200.140000 6.380000 ;
      RECT 0.000000 4.180000 4.340000 6.380000 ;
      RECT 0.000000 1.130000 1200.140000 4.180000 ;
      RECT 1.100000 1.100000 1200.140000 1.130000 ;
      RECT 1.850000 0.000000 1199.460000 1.100000 ;
      RECT 0.000000 0.000000 0.950000 0.230000 ;
    LAYER met4 ;
      RECT 0.000000 926.060000 1200.140000 930.580000 ;
      RECT 6.540000 922.860000 1193.600000 926.060000 ;
      RECT 1192.600000 7.380000 1193.600000 922.860000 ;
      RECT 9.740000 7.380000 1190.400000 922.860000 ;
      RECT 6.540000 7.380000 7.540000 922.860000 ;
      RECT 1195.800000 4.180000 1200.140000 926.060000 ;
      RECT 6.540000 4.180000 1193.600000 7.380000 ;
      RECT 0.000000 4.180000 4.340000 926.060000 ;
      RECT 0.000000 0.000000 1200.140000 4.180000 ;
      RECT 0.000000 0.000000 1200.140000 930.580000 ;
  END
END soc_now_caravel_top

END LIBRARY
