VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO soc_now_caravel_top
  CLASS BLOCK ;
  FOREIGN soc_now_caravel_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 1082.420 BY 1093.140 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 1089.140 728.090 1093.140 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1013.240 1082.420 1013.840 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 408.040 1082.420 408.640 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 1089.140 808.590 1093.140 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 197.240 1082.420 197.840 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 6.840 1082.420 7.440 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 901.040 1082.420 901.640 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 1089.140 634.710 1093.140 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 295.840 1082.420 296.440 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 1089.140 734.530 1093.140 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 1089.140 966.370 1093.140 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 982.640 1082.420 983.240 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1088.040 1082.420 1088.640 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 1089.140 380.330 1093.140 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 1089.140 509.130 1093.140 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 217.640 1082.420 218.240 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 894.240 1082.420 894.840 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 921.440 1082.420 922.040 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 428.440 1082.420 429.040 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 1089.140 860.110 1093.140 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1089.140 299.830 1093.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1089.140 315.930 1093.140 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 1089.140 87.310 1093.140 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 1089.140 354.570 1093.140 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 1089.140 361.010 1093.140 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1089.140 48.670 1093.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 850.040 1082.420 850.640 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 238.040 1082.420 238.640 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 1089.140 534.890 1093.140 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 112.240 1082.420 112.840 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 1089.140 1053.310 1093.140 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 204.040 1082.420 204.640 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 1089.140 1059.750 1093.140 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1089.140 167.810 1093.140 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 289.040 1082.420 289.640 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1089.140 0.370 1093.140 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 1089.140 740.970 1093.140 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 1089.140 406.090 1093.140 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 173.440 1082.420 174.040 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 1089.140 940.610 1093.140 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1081.240 1082.420 1081.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 1089.140 1027.550 1093.140 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 506.640 1082.420 507.240 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 870.440 1082.420 871.040 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 47.640 1082.420 48.240 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 1089.140 106.630 1093.140 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 1089.140 1008.230 1093.140 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 822.840 1082.420 823.440 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 462.440 1082.420 463.040 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 1089.140 187.130 1093.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 975.840 1082.420 976.440 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 1089.140 979.250 1093.140 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 139.440 1082.420 140.040 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 1089.140 567.090 1093.140 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 1089.140 228.990 1093.140 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 1089.140 74.430 1093.140 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 907.840 1082.420 908.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 1089.140 786.050 1093.140 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 1089.140 499.470 1093.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 1089.140 13.250 1093.140 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 771.840 1082.420 772.440 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 1089.140 866.550 1093.140 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 567.840 1082.420 568.440 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1089.140 113.070 1093.140 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 765.040 1082.420 765.640 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1089.140 399.650 1093.140 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 1089.140 554.210 1093.140 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 1089.140 335.250 1093.140 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 190.440 1082.420 191.040 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 744.640 1082.420 745.240 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 724.240 1082.420 724.840 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 493.040 1082.420 493.640 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 1089.140 879.430 1093.140 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 1089.140 766.730 1093.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 690.240 1082.420 690.840 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 343.440 1082.420 344.040 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 1089.140 341.690 1093.140 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 1089.140 473.710 1093.140 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 1089.140 328.810 1093.140 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1026.840 1082.420 1027.440 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 442.040 1082.420 442.640 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1089.140 19.690 1093.140 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 1089.140 306.270 1093.140 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 1089.140 61.550 1093.140 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 1089.140 628.270 1093.140 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1040.440 1082.420 1041.040 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 469.240 1082.420 469.840 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 717.440 1082.420 718.040 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1089.140 454.390 1093.140 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 809.240 1082.420 809.840 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 1089.140 422.190 1093.140 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 697.040 1082.420 697.640 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 435.240 1082.420 435.840 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 1089.140 821.470 1093.140 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 105.440 1082.420 106.040 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 731.040 1082.420 731.640 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 1089.140 934.170 1093.140 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 1089.140 393.210 1093.140 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 843.240 1082.420 843.840 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 0.040 1082.420 0.640 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 1089.140 621.830 1093.140 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.040 4.000 935.640 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 119.040 1082.420 119.640 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1089.140 67.990 1093.140 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 1089.140 435.070 1093.140 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 533.840 1082.420 534.440 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 1089.140 241.870 1093.140 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1089.140 560.650 1093.140 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 316.240 1082.420 316.840 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1089.140 100.190 1093.140 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 554.240 1082.420 554.840 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 1089.140 441.510 1093.140 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 1089.140 267.630 1093.140 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 357.040 1082.420 357.640 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 605.240 1082.420 605.840 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 639.240 1082.420 639.840 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 1089.140 174.250 1093.140 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 1089.140 1066.190 1093.140 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 710.640 1082.420 711.240 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 969.040 1082.420 969.640 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 598.440 1082.420 599.040 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 1089.140 673.350 1093.140 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 680.040 1082.420 680.640 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 547.440 1082.420 548.040 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 1089.140 708.770 1093.140 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 1089.140 1021.110 1093.140 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 336.640 1082.420 337.240 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 877.240 1082.420 877.840 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 941.840 1082.420 942.440 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 1089.140 834.350 1093.140 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 377.440 1082.420 378.040 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 1089.140 322.370 1093.140 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 98.640 1082.420 99.240 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 1089.140 927.730 1093.140 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 856.840 1082.420 857.440 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 414.840 1082.420 415.440 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 1089.140 985.690 1093.140 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 1089.140 386.770 1093.140 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 591.640 1082.420 592.240 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 1089.140 815.030 1093.140 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 1089.140 348.130 1093.140 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 1089.140 679.790 1093.140 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 829.640 1082.420 830.240 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 1089.140 486.590 1093.140 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 999.640 1082.420 1000.240 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 1089.140 760.290 1093.140 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 520.240 1082.420 520.840 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 1089.140 660.470 1093.140 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 625.640 1082.420 626.240 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 272.040 1082.420 272.640 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 1089.140 953.490 1093.140 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 166.640 1082.420 167.240 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 499.840 1082.420 500.440 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 703.840 1082.420 704.440 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 1089.140 802.150 1093.140 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 231.240 1082.420 231.840 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 1089.140 93.750 1093.140 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 159.840 1082.420 160.440 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1089.140 129.170 1093.140 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 513.440 1082.420 514.040 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 323.040 1082.420 323.640 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 989.440 1082.420 990.040 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 1089.140 1001.790 1093.140 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1089.140 35.790 1093.140 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 1089.140 222.550 1093.140 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 1089.140 193.570 1093.140 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 652.840 1082.420 653.440 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 574.640 1082.420 575.240 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 1089.140 206.450 1093.140 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 20.440 1082.420 21.040 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 1089.140 592.850 1093.140 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 244.840 1082.420 245.440 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 251.640 1082.420 252.240 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 1089.140 959.930 1093.140 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 1089.140 248.310 1093.140 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 1089.140 579.970 1093.140 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 1089.140 686.230 1093.140 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 125.840 1082.420 126.440 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1089.140 180.690 1093.140 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 91.840 1082.420 92.440 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 1089.140 415.750 1093.140 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 448.840 1082.420 449.440 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 1089.140 55.110 1093.140 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 1089.140 274.070 1093.140 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 1089.140 586.410 1093.140 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 1089.140 6.810 1093.140 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 1089.140 972.810 1093.140 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 1089.140 753.850 1093.140 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1089.140 428.630 1093.140 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 1089.140 161.370 1093.140 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 1089.140 921.290 1093.140 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 1089.140 885.870 1093.140 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 646.040 1082.420 646.640 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 282.240 1082.420 282.840 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 1089.140 261.190 1093.140 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 1089.140 148.490 1093.140 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 265.240 1082.420 265.840 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 1089.140 280.510 1093.140 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 1089.140 1014.670 1093.140 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1060.840 1082.420 1061.440 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 13.640 1082.420 14.240 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 618.840 1082.420 619.440 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 1089.140 367.450 1093.140 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 1089.140 493.030 1093.140 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 0.000 930.950 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 1089.140 547.770 1093.140 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1089.140 1072.630 1093.140 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 1089.140 853.670 1093.140 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 1089.140 827.910 1093.140 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 27.240 1082.420 27.840 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 1089.140 29.350 1093.140 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 1089.140 1040.430 1093.140 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 153.040 1082.420 153.640 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 1089.140 847.230 1093.140 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 1089.140 995.350 1093.140 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1089.140 779.610 1093.140 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 884.040 1082.420 884.640 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 612.040 1082.420 612.640 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 1089.140 573.530 1093.140 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 455.640 1082.420 456.240 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1089.140 80.870 1093.140 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 659.640 1082.420 660.240 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1089.140 212.890 1093.140 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 1089.140 615.390 1093.140 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 394.440 1082.420 395.040 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 561.040 1082.420 561.640 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 302.640 1082.420 303.240 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 795.640 1082.420 796.240 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 1089.140 608.950 1093.140 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 210.840 1082.420 211.440 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 183.640 1082.420 184.240 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1067.640 1082.420 1068.240 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 486.240 1082.420 486.840 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 401.240 1082.420 401.840 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 1089.140 901.970 1093.140 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 632.440 1082.420 633.040 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 1089.140 1033.990 1093.140 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 1089.140 1046.870 1093.140 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 85.040 1082.420 85.640 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1089.140 480.150 1093.140 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1033.640 1082.420 1034.240 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 0.000 966.370 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 0.000 1037.210 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 350.240 1082.420 350.840 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 935.040 1082.420 935.640 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 1089.140 515.570 1093.140 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 1089.140 467.270 1093.140 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1047.240 1082.420 1047.840 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1089.140 235.430 1093.140 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 914.640 1082.420 915.240 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 1089.140 647.590 1093.140 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 1089.140 840.790 1093.140 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 1089.140 895.530 1093.140 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 1089.140 908.410 1093.140 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 1089.140 541.330 1093.140 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 224.440 1082.420 225.040 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 1089.140 522.010 1093.140 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 785.440 1082.420 786.040 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1020.040 1082.420 1020.640 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 132.640 1082.420 133.240 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 962.240 1082.420 962.840 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 1089.140 373.890 1093.140 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 802.440 1082.420 803.040 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 0.000 924.510 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 1089.140 641.150 1093.140 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 258.440 1082.420 259.040 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 1089.140 293.390 1093.140 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 34.040 1082.420 34.640 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 758.240 1082.420 758.840 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 948.640 1082.420 949.240 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 54.440 1082.420 55.040 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 1089.140 42.230 1093.140 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 1087.440 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 1084.460 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 1085.840 1084.460 1087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1082.860 3.280 1084.460 1087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.720 -0.020 26.320 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.720 -0.020 206.320 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.720 457.180 206.320 490.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.720 907.180 206.320 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.720 -0.020 386.320 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.720 457.800 386.320 490.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.720 907.800 386.320 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 564.720 -0.020 566.320 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 744.720 -0.020 746.320 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 924.720 -0.020 926.320 1090.740 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 30.080 1087.760 31.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 210.080 1087.760 211.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 390.080 1087.760 391.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 570.080 1087.760 571.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 750.080 1087.760 751.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 930.080 1087.760 931.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 24.720 470.100 569.620 471.700 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 1090.740 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 1087.760 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1089.140 1087.760 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 1086.160 -0.020 1087.760 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.020 -0.020 29.620 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.020 -0.020 209.620 39.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.020 457.800 209.620 489.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.020 907.800 209.620 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 388.020 -0.020 389.620 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 388.020 457.180 389.620 490.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 388.020 907.180 389.620 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.020 -0.020 569.620 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 748.020 -0.020 749.620 1090.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 928.020 -0.020 929.620 1090.740 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 33.380 1087.760 34.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 213.380 1087.760 214.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 393.380 1087.760 394.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 573.380 1087.760 574.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 753.380 1087.760 754.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 933.380 1087.760 934.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 24.720 473.500 569.620 475.100 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 329.840 1082.420 330.440 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 540.640 1082.420 541.240 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 1089.140 447.950 1093.140 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 1089.140 200.010 1093.140 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1006.440 1082.420 1007.040 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 928.240 1082.420 928.840 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 836.440 1082.420 837.040 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 476.040 1082.420 476.640 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 40.840 1082.420 41.440 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1089.140 460.830 1093.140 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 363.840 1082.420 364.440 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1089.140 135.610 1093.140 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 778.640 1082.420 779.240 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 1089.140 947.050 1093.140 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 1089.140 666.910 1093.140 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 581.440 1082.420 582.040 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1089.140 654.030 1093.140 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 61.240 1082.420 61.840 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 387.640 1082.420 388.240 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 1089.140 154.930 1093.140 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 1089.140 1079.070 1093.140 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 666.440 1082.420 667.040 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 1089.140 599.290 1093.140 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 1089.140 872.990 1093.140 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 982.640 4.000 983.240 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 751.440 1082.420 752.040 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 1089.140 914.850 1093.140 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 955.440 1082.420 956.040 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 421.640 1082.420 422.240 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 1089.140 792.490 1093.140 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 1089.140 142.050 1093.140 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 737.840 1082.420 738.440 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 370.640 1082.420 371.240 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 68.040 1082.420 68.640 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 1089.140 773.170 1093.140 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1054.040 1082.420 1054.640 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 78.240 1082.420 78.840 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 673.240 1082.420 673.840 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 1074.440 1082.420 1075.040 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 1089.140 747.410 1093.140 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 146.240 1082.420 146.840 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 1089.140 715.210 1093.140 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 1089.140 254.750 1093.140 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 1089.140 528.450 1093.140 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 1089.140 286.950 1093.140 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1089.140 721.650 1093.140 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 309.440 1082.420 310.040 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 863.640 1082.420 864.240 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 816.040 1082.420 816.640 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 1089.140 702.330 1093.140 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 1089.140 692.670 1093.140 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1089.140 122.730 1093.140 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1078.420 527.040 1082.420 527.640 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 7.905 1082.235 1081.455 ;
      LAYER met1 ;
        RECT 0.070 1.400 1082.310 1081.500 ;
      LAYER met2 ;
        RECT 0.650 1088.860 6.250 1089.770 ;
        RECT 7.090 1088.860 12.690 1089.770 ;
        RECT 13.530 1088.860 19.130 1089.770 ;
        RECT 19.970 1088.860 28.790 1089.770 ;
        RECT 29.630 1088.860 35.230 1089.770 ;
        RECT 36.070 1088.860 41.670 1089.770 ;
        RECT 42.510 1088.860 48.110 1089.770 ;
        RECT 48.950 1088.860 54.550 1089.770 ;
        RECT 55.390 1088.860 60.990 1089.770 ;
        RECT 61.830 1088.860 67.430 1089.770 ;
        RECT 68.270 1088.860 73.870 1089.770 ;
        RECT 74.710 1088.860 80.310 1089.770 ;
        RECT 81.150 1088.860 86.750 1089.770 ;
        RECT 87.590 1088.860 93.190 1089.770 ;
        RECT 94.030 1088.860 99.630 1089.770 ;
        RECT 100.470 1088.860 106.070 1089.770 ;
        RECT 106.910 1088.860 112.510 1089.770 ;
        RECT 113.350 1088.860 122.170 1089.770 ;
        RECT 123.010 1088.860 128.610 1089.770 ;
        RECT 129.450 1088.860 135.050 1089.770 ;
        RECT 135.890 1088.860 141.490 1089.770 ;
        RECT 142.330 1088.860 147.930 1089.770 ;
        RECT 148.770 1088.860 154.370 1089.770 ;
        RECT 155.210 1088.860 160.810 1089.770 ;
        RECT 161.650 1088.860 167.250 1089.770 ;
        RECT 168.090 1088.860 173.690 1089.770 ;
        RECT 174.530 1088.860 180.130 1089.770 ;
        RECT 180.970 1088.860 186.570 1089.770 ;
        RECT 187.410 1088.860 193.010 1089.770 ;
        RECT 193.850 1088.860 199.450 1089.770 ;
        RECT 200.290 1088.860 205.890 1089.770 ;
        RECT 206.730 1088.860 212.330 1089.770 ;
        RECT 213.170 1088.860 221.990 1089.770 ;
        RECT 222.830 1088.860 228.430 1089.770 ;
        RECT 229.270 1088.860 234.870 1089.770 ;
        RECT 235.710 1088.860 241.310 1089.770 ;
        RECT 242.150 1088.860 247.750 1089.770 ;
        RECT 248.590 1088.860 254.190 1089.770 ;
        RECT 255.030 1088.860 260.630 1089.770 ;
        RECT 261.470 1088.860 267.070 1089.770 ;
        RECT 267.910 1088.860 273.510 1089.770 ;
        RECT 274.350 1088.860 279.950 1089.770 ;
        RECT 280.790 1088.860 286.390 1089.770 ;
        RECT 287.230 1088.860 292.830 1089.770 ;
        RECT 293.670 1088.860 299.270 1089.770 ;
        RECT 300.110 1088.860 305.710 1089.770 ;
        RECT 306.550 1088.860 315.370 1089.770 ;
        RECT 316.210 1088.860 321.810 1089.770 ;
        RECT 322.650 1088.860 328.250 1089.770 ;
        RECT 329.090 1088.860 334.690 1089.770 ;
        RECT 335.530 1088.860 341.130 1089.770 ;
        RECT 341.970 1088.860 347.570 1089.770 ;
        RECT 348.410 1088.860 354.010 1089.770 ;
        RECT 354.850 1088.860 360.450 1089.770 ;
        RECT 361.290 1088.860 366.890 1089.770 ;
        RECT 367.730 1088.860 373.330 1089.770 ;
        RECT 374.170 1088.860 379.770 1089.770 ;
        RECT 380.610 1088.860 386.210 1089.770 ;
        RECT 387.050 1088.860 392.650 1089.770 ;
        RECT 393.490 1088.860 399.090 1089.770 ;
        RECT 399.930 1088.860 405.530 1089.770 ;
        RECT 406.370 1088.860 415.190 1089.770 ;
        RECT 416.030 1088.860 421.630 1089.770 ;
        RECT 422.470 1088.860 428.070 1089.770 ;
        RECT 428.910 1088.860 434.510 1089.770 ;
        RECT 435.350 1088.860 440.950 1089.770 ;
        RECT 441.790 1088.860 447.390 1089.770 ;
        RECT 448.230 1088.860 453.830 1089.770 ;
        RECT 454.670 1088.860 460.270 1089.770 ;
        RECT 461.110 1088.860 466.710 1089.770 ;
        RECT 467.550 1088.860 473.150 1089.770 ;
        RECT 473.990 1088.860 479.590 1089.770 ;
        RECT 480.430 1088.860 486.030 1089.770 ;
        RECT 486.870 1088.860 492.470 1089.770 ;
        RECT 493.310 1088.860 498.910 1089.770 ;
        RECT 499.750 1088.860 508.570 1089.770 ;
        RECT 509.410 1088.860 515.010 1089.770 ;
        RECT 515.850 1088.860 521.450 1089.770 ;
        RECT 522.290 1088.860 527.890 1089.770 ;
        RECT 528.730 1088.860 534.330 1089.770 ;
        RECT 535.170 1088.860 540.770 1089.770 ;
        RECT 541.610 1088.860 547.210 1089.770 ;
        RECT 548.050 1088.860 553.650 1089.770 ;
        RECT 554.490 1088.860 560.090 1089.770 ;
        RECT 560.930 1088.860 566.530 1089.770 ;
        RECT 567.370 1088.860 572.970 1089.770 ;
        RECT 573.810 1088.860 579.410 1089.770 ;
        RECT 580.250 1088.860 585.850 1089.770 ;
        RECT 586.690 1088.860 592.290 1089.770 ;
        RECT 593.130 1088.860 598.730 1089.770 ;
        RECT 599.570 1088.860 608.390 1089.770 ;
        RECT 609.230 1088.860 614.830 1089.770 ;
        RECT 615.670 1088.860 621.270 1089.770 ;
        RECT 622.110 1088.860 627.710 1089.770 ;
        RECT 628.550 1088.860 634.150 1089.770 ;
        RECT 634.990 1088.860 640.590 1089.770 ;
        RECT 641.430 1088.860 647.030 1089.770 ;
        RECT 647.870 1088.860 653.470 1089.770 ;
        RECT 654.310 1088.860 659.910 1089.770 ;
        RECT 660.750 1088.860 666.350 1089.770 ;
        RECT 667.190 1088.860 672.790 1089.770 ;
        RECT 673.630 1088.860 679.230 1089.770 ;
        RECT 680.070 1088.860 685.670 1089.770 ;
        RECT 686.510 1088.860 692.110 1089.770 ;
        RECT 692.950 1088.860 701.770 1089.770 ;
        RECT 702.610 1088.860 708.210 1089.770 ;
        RECT 709.050 1088.860 714.650 1089.770 ;
        RECT 715.490 1088.860 721.090 1089.770 ;
        RECT 721.930 1088.860 727.530 1089.770 ;
        RECT 728.370 1088.860 733.970 1089.770 ;
        RECT 734.810 1088.860 740.410 1089.770 ;
        RECT 741.250 1088.860 746.850 1089.770 ;
        RECT 747.690 1088.860 753.290 1089.770 ;
        RECT 754.130 1088.860 759.730 1089.770 ;
        RECT 760.570 1088.860 766.170 1089.770 ;
        RECT 767.010 1088.860 772.610 1089.770 ;
        RECT 773.450 1088.860 779.050 1089.770 ;
        RECT 779.890 1088.860 785.490 1089.770 ;
        RECT 786.330 1088.860 791.930 1089.770 ;
        RECT 792.770 1088.860 801.590 1089.770 ;
        RECT 802.430 1088.860 808.030 1089.770 ;
        RECT 808.870 1088.860 814.470 1089.770 ;
        RECT 815.310 1088.860 820.910 1089.770 ;
        RECT 821.750 1088.860 827.350 1089.770 ;
        RECT 828.190 1088.860 833.790 1089.770 ;
        RECT 834.630 1088.860 840.230 1089.770 ;
        RECT 841.070 1088.860 846.670 1089.770 ;
        RECT 847.510 1088.860 853.110 1089.770 ;
        RECT 853.950 1088.860 859.550 1089.770 ;
        RECT 860.390 1088.860 865.990 1089.770 ;
        RECT 866.830 1088.860 872.430 1089.770 ;
        RECT 873.270 1088.860 878.870 1089.770 ;
        RECT 879.710 1088.860 885.310 1089.770 ;
        RECT 886.150 1088.860 894.970 1089.770 ;
        RECT 895.810 1088.860 901.410 1089.770 ;
        RECT 902.250 1088.860 907.850 1089.770 ;
        RECT 908.690 1088.860 914.290 1089.770 ;
        RECT 915.130 1088.860 920.730 1089.770 ;
        RECT 921.570 1088.860 927.170 1089.770 ;
        RECT 928.010 1088.860 933.610 1089.770 ;
        RECT 934.450 1088.860 940.050 1089.770 ;
        RECT 940.890 1088.860 946.490 1089.770 ;
        RECT 947.330 1088.860 952.930 1089.770 ;
        RECT 953.770 1088.860 959.370 1089.770 ;
        RECT 960.210 1088.860 965.810 1089.770 ;
        RECT 966.650 1088.860 972.250 1089.770 ;
        RECT 973.090 1088.860 978.690 1089.770 ;
        RECT 979.530 1088.860 985.130 1089.770 ;
        RECT 985.970 1088.860 994.790 1089.770 ;
        RECT 995.630 1088.860 1001.230 1089.770 ;
        RECT 1002.070 1088.860 1007.670 1089.770 ;
        RECT 1008.510 1088.860 1014.110 1089.770 ;
        RECT 1014.950 1088.860 1020.550 1089.770 ;
        RECT 1021.390 1088.860 1026.990 1089.770 ;
        RECT 1027.830 1088.860 1033.430 1089.770 ;
        RECT 1034.270 1088.860 1039.870 1089.770 ;
        RECT 1040.710 1088.860 1046.310 1089.770 ;
        RECT 1047.150 1088.860 1052.750 1089.770 ;
        RECT 1053.590 1088.860 1059.190 1089.770 ;
        RECT 1060.030 1088.860 1065.630 1089.770 ;
        RECT 1066.470 1088.860 1072.070 1089.770 ;
        RECT 1072.910 1088.860 1078.510 1089.770 ;
        RECT 1079.350 1088.860 1082.280 1089.770 ;
        RECT 0.100 4.280 1082.280 1088.860 ;
        RECT 0.650 1.370 6.250 4.280 ;
        RECT 7.090 1.370 12.690 4.280 ;
        RECT 13.530 1.370 19.130 4.280 ;
        RECT 19.970 1.370 25.570 4.280 ;
        RECT 26.410 1.370 32.010 4.280 ;
        RECT 32.850 1.370 38.450 4.280 ;
        RECT 39.290 1.370 44.890 4.280 ;
        RECT 45.730 1.370 51.330 4.280 ;
        RECT 52.170 1.370 57.770 4.280 ;
        RECT 58.610 1.370 64.210 4.280 ;
        RECT 65.050 1.370 70.650 4.280 ;
        RECT 71.490 1.370 77.090 4.280 ;
        RECT 77.930 1.370 83.530 4.280 ;
        RECT 84.370 1.370 89.970 4.280 ;
        RECT 90.810 1.370 99.630 4.280 ;
        RECT 100.470 1.370 106.070 4.280 ;
        RECT 106.910 1.370 112.510 4.280 ;
        RECT 113.350 1.370 118.950 4.280 ;
        RECT 119.790 1.370 125.390 4.280 ;
        RECT 126.230 1.370 131.830 4.280 ;
        RECT 132.670 1.370 138.270 4.280 ;
        RECT 139.110 1.370 144.710 4.280 ;
        RECT 145.550 1.370 151.150 4.280 ;
        RECT 151.990 1.370 157.590 4.280 ;
        RECT 158.430 1.370 164.030 4.280 ;
        RECT 164.870 1.370 170.470 4.280 ;
        RECT 171.310 1.370 176.910 4.280 ;
        RECT 177.750 1.370 183.350 4.280 ;
        RECT 184.190 1.370 193.010 4.280 ;
        RECT 193.850 1.370 199.450 4.280 ;
        RECT 200.290 1.370 205.890 4.280 ;
        RECT 206.730 1.370 212.330 4.280 ;
        RECT 213.170 1.370 218.770 4.280 ;
        RECT 219.610 1.370 225.210 4.280 ;
        RECT 226.050 1.370 231.650 4.280 ;
        RECT 232.490 1.370 238.090 4.280 ;
        RECT 238.930 1.370 244.530 4.280 ;
        RECT 245.370 1.370 250.970 4.280 ;
        RECT 251.810 1.370 257.410 4.280 ;
        RECT 258.250 1.370 263.850 4.280 ;
        RECT 264.690 1.370 270.290 4.280 ;
        RECT 271.130 1.370 276.730 4.280 ;
        RECT 277.570 1.370 283.170 4.280 ;
        RECT 284.010 1.370 292.830 4.280 ;
        RECT 293.670 1.370 299.270 4.280 ;
        RECT 300.110 1.370 305.710 4.280 ;
        RECT 306.550 1.370 312.150 4.280 ;
        RECT 312.990 1.370 318.590 4.280 ;
        RECT 319.430 1.370 325.030 4.280 ;
        RECT 325.870 1.370 331.470 4.280 ;
        RECT 332.310 1.370 337.910 4.280 ;
        RECT 338.750 1.370 344.350 4.280 ;
        RECT 345.190 1.370 350.790 4.280 ;
        RECT 351.630 1.370 357.230 4.280 ;
        RECT 358.070 1.370 363.670 4.280 ;
        RECT 364.510 1.370 370.110 4.280 ;
        RECT 370.950 1.370 376.550 4.280 ;
        RECT 377.390 1.370 386.210 4.280 ;
        RECT 387.050 1.370 392.650 4.280 ;
        RECT 393.490 1.370 399.090 4.280 ;
        RECT 399.930 1.370 405.530 4.280 ;
        RECT 406.370 1.370 411.970 4.280 ;
        RECT 412.810 1.370 418.410 4.280 ;
        RECT 419.250 1.370 424.850 4.280 ;
        RECT 425.690 1.370 431.290 4.280 ;
        RECT 432.130 1.370 437.730 4.280 ;
        RECT 438.570 1.370 444.170 4.280 ;
        RECT 445.010 1.370 450.610 4.280 ;
        RECT 451.450 1.370 457.050 4.280 ;
        RECT 457.890 1.370 463.490 4.280 ;
        RECT 464.330 1.370 469.930 4.280 ;
        RECT 470.770 1.370 476.370 4.280 ;
        RECT 477.210 1.370 486.030 4.280 ;
        RECT 486.870 1.370 492.470 4.280 ;
        RECT 493.310 1.370 498.910 4.280 ;
        RECT 499.750 1.370 505.350 4.280 ;
        RECT 506.190 1.370 511.790 4.280 ;
        RECT 512.630 1.370 518.230 4.280 ;
        RECT 519.070 1.370 524.670 4.280 ;
        RECT 525.510 1.370 531.110 4.280 ;
        RECT 531.950 1.370 537.550 4.280 ;
        RECT 538.390 1.370 543.990 4.280 ;
        RECT 544.830 1.370 550.430 4.280 ;
        RECT 551.270 1.370 556.870 4.280 ;
        RECT 557.710 1.370 563.310 4.280 ;
        RECT 564.150 1.370 569.750 4.280 ;
        RECT 570.590 1.370 579.410 4.280 ;
        RECT 580.250 1.370 585.850 4.280 ;
        RECT 586.690 1.370 592.290 4.280 ;
        RECT 593.130 1.370 598.730 4.280 ;
        RECT 599.570 1.370 605.170 4.280 ;
        RECT 606.010 1.370 611.610 4.280 ;
        RECT 612.450 1.370 618.050 4.280 ;
        RECT 618.890 1.370 624.490 4.280 ;
        RECT 625.330 1.370 630.930 4.280 ;
        RECT 631.770 1.370 637.370 4.280 ;
        RECT 638.210 1.370 643.810 4.280 ;
        RECT 644.650 1.370 650.250 4.280 ;
        RECT 651.090 1.370 656.690 4.280 ;
        RECT 657.530 1.370 663.130 4.280 ;
        RECT 663.970 1.370 669.570 4.280 ;
        RECT 670.410 1.370 679.230 4.280 ;
        RECT 680.070 1.370 685.670 4.280 ;
        RECT 686.510 1.370 692.110 4.280 ;
        RECT 692.950 1.370 698.550 4.280 ;
        RECT 699.390 1.370 704.990 4.280 ;
        RECT 705.830 1.370 711.430 4.280 ;
        RECT 712.270 1.370 717.870 4.280 ;
        RECT 718.710 1.370 724.310 4.280 ;
        RECT 725.150 1.370 730.750 4.280 ;
        RECT 731.590 1.370 737.190 4.280 ;
        RECT 738.030 1.370 743.630 4.280 ;
        RECT 744.470 1.370 750.070 4.280 ;
        RECT 750.910 1.370 756.510 4.280 ;
        RECT 757.350 1.370 762.950 4.280 ;
        RECT 763.790 1.370 772.610 4.280 ;
        RECT 773.450 1.370 779.050 4.280 ;
        RECT 779.890 1.370 785.490 4.280 ;
        RECT 786.330 1.370 791.930 4.280 ;
        RECT 792.770 1.370 798.370 4.280 ;
        RECT 799.210 1.370 804.810 4.280 ;
        RECT 805.650 1.370 811.250 4.280 ;
        RECT 812.090 1.370 817.690 4.280 ;
        RECT 818.530 1.370 824.130 4.280 ;
        RECT 824.970 1.370 830.570 4.280 ;
        RECT 831.410 1.370 837.010 4.280 ;
        RECT 837.850 1.370 843.450 4.280 ;
        RECT 844.290 1.370 849.890 4.280 ;
        RECT 850.730 1.370 856.330 4.280 ;
        RECT 857.170 1.370 862.770 4.280 ;
        RECT 863.610 1.370 872.430 4.280 ;
        RECT 873.270 1.370 878.870 4.280 ;
        RECT 879.710 1.370 885.310 4.280 ;
        RECT 886.150 1.370 891.750 4.280 ;
        RECT 892.590 1.370 898.190 4.280 ;
        RECT 899.030 1.370 904.630 4.280 ;
        RECT 905.470 1.370 911.070 4.280 ;
        RECT 911.910 1.370 917.510 4.280 ;
        RECT 918.350 1.370 923.950 4.280 ;
        RECT 924.790 1.370 930.390 4.280 ;
        RECT 931.230 1.370 936.830 4.280 ;
        RECT 937.670 1.370 943.270 4.280 ;
        RECT 944.110 1.370 949.710 4.280 ;
        RECT 950.550 1.370 956.150 4.280 ;
        RECT 956.990 1.370 965.810 4.280 ;
        RECT 966.650 1.370 972.250 4.280 ;
        RECT 973.090 1.370 978.690 4.280 ;
        RECT 979.530 1.370 985.130 4.280 ;
        RECT 985.970 1.370 991.570 4.280 ;
        RECT 992.410 1.370 998.010 4.280 ;
        RECT 998.850 1.370 1004.450 4.280 ;
        RECT 1005.290 1.370 1010.890 4.280 ;
        RECT 1011.730 1.370 1017.330 4.280 ;
        RECT 1018.170 1.370 1023.770 4.280 ;
        RECT 1024.610 1.370 1030.210 4.280 ;
        RECT 1031.050 1.370 1036.650 4.280 ;
        RECT 1037.490 1.370 1043.090 4.280 ;
        RECT 1043.930 1.370 1049.530 4.280 ;
        RECT 1050.370 1.370 1055.970 4.280 ;
        RECT 1056.810 1.370 1065.630 4.280 ;
        RECT 1066.470 1.370 1072.070 4.280 ;
        RECT 1072.910 1.370 1078.510 4.280 ;
        RECT 1079.350 1.370 1082.280 4.280 ;
      LAYER met3 ;
        RECT 4.400 1080.840 1078.020 1081.705 ;
        RECT 4.000 1075.440 1078.420 1080.840 ;
        RECT 4.400 1074.040 1078.020 1075.440 ;
        RECT 4.000 1068.640 1078.420 1074.040 ;
        RECT 4.400 1067.240 1078.020 1068.640 ;
        RECT 4.000 1061.840 1078.420 1067.240 ;
        RECT 4.400 1060.440 1078.020 1061.840 ;
        RECT 4.000 1055.040 1078.420 1060.440 ;
        RECT 4.400 1053.640 1078.020 1055.040 ;
        RECT 4.000 1048.240 1078.420 1053.640 ;
        RECT 4.400 1046.840 1078.020 1048.240 ;
        RECT 4.000 1041.440 1078.420 1046.840 ;
        RECT 4.400 1040.040 1078.020 1041.440 ;
        RECT 4.000 1034.640 1078.420 1040.040 ;
        RECT 4.400 1033.240 1078.020 1034.640 ;
        RECT 4.000 1027.840 1078.420 1033.240 ;
        RECT 4.400 1026.440 1078.020 1027.840 ;
        RECT 4.000 1021.040 1078.420 1026.440 ;
        RECT 4.400 1019.640 1078.020 1021.040 ;
        RECT 4.000 1014.240 1078.420 1019.640 ;
        RECT 4.000 1012.840 1078.020 1014.240 ;
        RECT 4.000 1010.840 1078.420 1012.840 ;
        RECT 4.400 1009.440 1078.420 1010.840 ;
        RECT 4.000 1007.440 1078.420 1009.440 ;
        RECT 4.000 1006.040 1078.020 1007.440 ;
        RECT 4.000 1004.040 1078.420 1006.040 ;
        RECT 4.400 1002.640 1078.420 1004.040 ;
        RECT 4.000 1000.640 1078.420 1002.640 ;
        RECT 4.000 999.240 1078.020 1000.640 ;
        RECT 4.000 997.240 1078.420 999.240 ;
        RECT 4.400 995.840 1078.420 997.240 ;
        RECT 4.000 990.440 1078.420 995.840 ;
        RECT 4.400 989.040 1078.020 990.440 ;
        RECT 4.000 983.640 1078.420 989.040 ;
        RECT 4.400 982.240 1078.020 983.640 ;
        RECT 4.000 976.840 1078.420 982.240 ;
        RECT 4.400 975.440 1078.020 976.840 ;
        RECT 4.000 970.040 1078.420 975.440 ;
        RECT 4.400 968.640 1078.020 970.040 ;
        RECT 4.000 963.240 1078.420 968.640 ;
        RECT 4.400 961.840 1078.020 963.240 ;
        RECT 4.000 956.440 1078.420 961.840 ;
        RECT 4.400 955.040 1078.020 956.440 ;
        RECT 4.000 949.640 1078.420 955.040 ;
        RECT 4.400 948.240 1078.020 949.640 ;
        RECT 4.000 942.840 1078.420 948.240 ;
        RECT 4.400 941.440 1078.020 942.840 ;
        RECT 4.000 936.040 1078.420 941.440 ;
        RECT 4.400 934.640 1078.020 936.040 ;
        RECT 4.000 929.240 1078.420 934.640 ;
        RECT 4.400 927.840 1078.020 929.240 ;
        RECT 4.000 922.440 1078.420 927.840 ;
        RECT 4.400 921.040 1078.020 922.440 ;
        RECT 4.000 915.640 1078.420 921.040 ;
        RECT 4.000 914.240 1078.020 915.640 ;
        RECT 4.000 912.240 1078.420 914.240 ;
        RECT 4.400 910.840 1078.420 912.240 ;
        RECT 4.000 908.840 1078.420 910.840 ;
        RECT 4.000 907.440 1078.020 908.840 ;
        RECT 4.000 905.440 1078.420 907.440 ;
        RECT 4.400 904.040 1078.420 905.440 ;
        RECT 4.000 902.040 1078.420 904.040 ;
        RECT 4.000 900.640 1078.020 902.040 ;
        RECT 4.000 898.640 1078.420 900.640 ;
        RECT 4.400 897.240 1078.420 898.640 ;
        RECT 4.000 895.240 1078.420 897.240 ;
        RECT 4.000 893.840 1078.020 895.240 ;
        RECT 4.000 891.840 1078.420 893.840 ;
        RECT 4.400 890.440 1078.420 891.840 ;
        RECT 4.000 885.040 1078.420 890.440 ;
        RECT 4.400 883.640 1078.020 885.040 ;
        RECT 4.000 878.240 1078.420 883.640 ;
        RECT 4.400 876.840 1078.020 878.240 ;
        RECT 4.000 871.440 1078.420 876.840 ;
        RECT 4.400 870.040 1078.020 871.440 ;
        RECT 4.000 864.640 1078.420 870.040 ;
        RECT 4.400 863.240 1078.020 864.640 ;
        RECT 4.000 857.840 1078.420 863.240 ;
        RECT 4.400 856.440 1078.020 857.840 ;
        RECT 4.000 851.040 1078.420 856.440 ;
        RECT 4.400 849.640 1078.020 851.040 ;
        RECT 4.000 844.240 1078.420 849.640 ;
        RECT 4.400 842.840 1078.020 844.240 ;
        RECT 4.000 837.440 1078.420 842.840 ;
        RECT 4.400 836.040 1078.020 837.440 ;
        RECT 4.000 830.640 1078.420 836.040 ;
        RECT 4.400 829.240 1078.020 830.640 ;
        RECT 4.000 823.840 1078.420 829.240 ;
        RECT 4.400 822.440 1078.020 823.840 ;
        RECT 4.000 817.040 1078.420 822.440 ;
        RECT 4.400 815.640 1078.020 817.040 ;
        RECT 4.000 810.240 1078.420 815.640 ;
        RECT 4.000 808.840 1078.020 810.240 ;
        RECT 4.000 806.840 1078.420 808.840 ;
        RECT 4.400 805.440 1078.420 806.840 ;
        RECT 4.000 803.440 1078.420 805.440 ;
        RECT 4.000 802.040 1078.020 803.440 ;
        RECT 4.000 800.040 1078.420 802.040 ;
        RECT 4.400 798.640 1078.420 800.040 ;
        RECT 4.000 796.640 1078.420 798.640 ;
        RECT 4.000 795.240 1078.020 796.640 ;
        RECT 4.000 793.240 1078.420 795.240 ;
        RECT 4.400 791.840 1078.420 793.240 ;
        RECT 4.000 786.440 1078.420 791.840 ;
        RECT 4.400 785.040 1078.020 786.440 ;
        RECT 4.000 779.640 1078.420 785.040 ;
        RECT 4.400 778.240 1078.020 779.640 ;
        RECT 4.000 772.840 1078.420 778.240 ;
        RECT 4.400 771.440 1078.020 772.840 ;
        RECT 4.000 766.040 1078.420 771.440 ;
        RECT 4.400 764.640 1078.020 766.040 ;
        RECT 4.000 759.240 1078.420 764.640 ;
        RECT 4.400 757.840 1078.020 759.240 ;
        RECT 4.000 752.440 1078.420 757.840 ;
        RECT 4.400 751.040 1078.020 752.440 ;
        RECT 4.000 745.640 1078.420 751.040 ;
        RECT 4.400 744.240 1078.020 745.640 ;
        RECT 4.000 738.840 1078.420 744.240 ;
        RECT 4.400 737.440 1078.020 738.840 ;
        RECT 4.000 732.040 1078.420 737.440 ;
        RECT 4.400 730.640 1078.020 732.040 ;
        RECT 4.000 725.240 1078.420 730.640 ;
        RECT 4.400 723.840 1078.020 725.240 ;
        RECT 4.000 718.440 1078.420 723.840 ;
        RECT 4.400 717.040 1078.020 718.440 ;
        RECT 4.000 711.640 1078.420 717.040 ;
        RECT 4.000 710.240 1078.020 711.640 ;
        RECT 4.000 708.240 1078.420 710.240 ;
        RECT 4.400 706.840 1078.420 708.240 ;
        RECT 4.000 704.840 1078.420 706.840 ;
        RECT 4.000 703.440 1078.020 704.840 ;
        RECT 4.000 701.440 1078.420 703.440 ;
        RECT 4.400 700.040 1078.420 701.440 ;
        RECT 4.000 698.040 1078.420 700.040 ;
        RECT 4.000 696.640 1078.020 698.040 ;
        RECT 4.000 694.640 1078.420 696.640 ;
        RECT 4.400 693.240 1078.420 694.640 ;
        RECT 4.000 691.240 1078.420 693.240 ;
        RECT 4.000 689.840 1078.020 691.240 ;
        RECT 4.000 687.840 1078.420 689.840 ;
        RECT 4.400 686.440 1078.420 687.840 ;
        RECT 4.000 681.040 1078.420 686.440 ;
        RECT 4.400 679.640 1078.020 681.040 ;
        RECT 4.000 674.240 1078.420 679.640 ;
        RECT 4.400 672.840 1078.020 674.240 ;
        RECT 4.000 667.440 1078.420 672.840 ;
        RECT 4.400 666.040 1078.020 667.440 ;
        RECT 4.000 660.640 1078.420 666.040 ;
        RECT 4.400 659.240 1078.020 660.640 ;
        RECT 4.000 653.840 1078.420 659.240 ;
        RECT 4.400 652.440 1078.020 653.840 ;
        RECT 4.000 647.040 1078.420 652.440 ;
        RECT 4.400 645.640 1078.020 647.040 ;
        RECT 4.000 640.240 1078.420 645.640 ;
        RECT 4.400 638.840 1078.020 640.240 ;
        RECT 4.000 633.440 1078.420 638.840 ;
        RECT 4.400 632.040 1078.020 633.440 ;
        RECT 4.000 626.640 1078.420 632.040 ;
        RECT 4.400 625.240 1078.020 626.640 ;
        RECT 4.000 619.840 1078.420 625.240 ;
        RECT 4.400 618.440 1078.020 619.840 ;
        RECT 4.000 613.040 1078.420 618.440 ;
        RECT 4.400 611.640 1078.020 613.040 ;
        RECT 4.000 606.240 1078.420 611.640 ;
        RECT 4.000 604.840 1078.020 606.240 ;
        RECT 4.000 602.840 1078.420 604.840 ;
        RECT 4.400 601.440 1078.420 602.840 ;
        RECT 4.000 599.440 1078.420 601.440 ;
        RECT 4.000 598.040 1078.020 599.440 ;
        RECT 4.000 596.040 1078.420 598.040 ;
        RECT 4.400 594.640 1078.420 596.040 ;
        RECT 4.000 592.640 1078.420 594.640 ;
        RECT 4.000 591.240 1078.020 592.640 ;
        RECT 4.000 589.240 1078.420 591.240 ;
        RECT 4.400 587.840 1078.420 589.240 ;
        RECT 4.000 582.440 1078.420 587.840 ;
        RECT 4.400 581.040 1078.020 582.440 ;
        RECT 4.000 575.640 1078.420 581.040 ;
        RECT 4.400 574.240 1078.020 575.640 ;
        RECT 4.000 568.840 1078.420 574.240 ;
        RECT 4.400 567.440 1078.020 568.840 ;
        RECT 4.000 562.040 1078.420 567.440 ;
        RECT 4.400 560.640 1078.020 562.040 ;
        RECT 4.000 555.240 1078.420 560.640 ;
        RECT 4.400 553.840 1078.020 555.240 ;
        RECT 4.000 548.440 1078.420 553.840 ;
        RECT 4.400 547.040 1078.020 548.440 ;
        RECT 4.000 541.640 1078.420 547.040 ;
        RECT 4.400 540.240 1078.020 541.640 ;
        RECT 4.000 534.840 1078.420 540.240 ;
        RECT 4.400 533.440 1078.020 534.840 ;
        RECT 4.000 528.040 1078.420 533.440 ;
        RECT 4.400 526.640 1078.020 528.040 ;
        RECT 4.000 521.240 1078.420 526.640 ;
        RECT 4.400 519.840 1078.020 521.240 ;
        RECT 4.000 514.440 1078.420 519.840 ;
        RECT 4.400 513.040 1078.020 514.440 ;
        RECT 4.000 507.640 1078.420 513.040 ;
        RECT 4.000 506.240 1078.020 507.640 ;
        RECT 4.000 504.240 1078.420 506.240 ;
        RECT 4.400 502.840 1078.420 504.240 ;
        RECT 4.000 500.840 1078.420 502.840 ;
        RECT 4.000 499.440 1078.020 500.840 ;
        RECT 4.000 497.440 1078.420 499.440 ;
        RECT 4.400 496.040 1078.420 497.440 ;
        RECT 4.000 494.040 1078.420 496.040 ;
        RECT 4.000 492.640 1078.020 494.040 ;
        RECT 4.000 490.640 1078.420 492.640 ;
        RECT 4.400 489.240 1078.420 490.640 ;
        RECT 4.000 487.240 1078.420 489.240 ;
        RECT 4.000 485.840 1078.020 487.240 ;
        RECT 4.000 483.840 1078.420 485.840 ;
        RECT 4.400 482.440 1078.420 483.840 ;
        RECT 4.000 477.040 1078.420 482.440 ;
        RECT 4.400 475.640 1078.020 477.040 ;
        RECT 4.000 470.240 1078.420 475.640 ;
        RECT 4.400 468.840 1078.020 470.240 ;
        RECT 4.000 463.440 1078.420 468.840 ;
        RECT 4.400 462.040 1078.020 463.440 ;
        RECT 4.000 456.640 1078.420 462.040 ;
        RECT 4.400 455.240 1078.020 456.640 ;
        RECT 4.000 449.840 1078.420 455.240 ;
        RECT 4.400 448.440 1078.020 449.840 ;
        RECT 4.000 443.040 1078.420 448.440 ;
        RECT 4.400 441.640 1078.020 443.040 ;
        RECT 4.000 436.240 1078.420 441.640 ;
        RECT 4.400 434.840 1078.020 436.240 ;
        RECT 4.000 429.440 1078.420 434.840 ;
        RECT 4.400 428.040 1078.020 429.440 ;
        RECT 4.000 422.640 1078.420 428.040 ;
        RECT 4.400 421.240 1078.020 422.640 ;
        RECT 4.000 415.840 1078.420 421.240 ;
        RECT 4.400 414.440 1078.020 415.840 ;
        RECT 4.000 409.040 1078.420 414.440 ;
        RECT 4.400 407.640 1078.020 409.040 ;
        RECT 4.000 402.240 1078.420 407.640 ;
        RECT 4.000 400.840 1078.020 402.240 ;
        RECT 4.000 398.840 1078.420 400.840 ;
        RECT 4.400 397.440 1078.420 398.840 ;
        RECT 4.000 395.440 1078.420 397.440 ;
        RECT 4.000 394.040 1078.020 395.440 ;
        RECT 4.000 392.040 1078.420 394.040 ;
        RECT 4.400 390.640 1078.420 392.040 ;
        RECT 4.000 388.640 1078.420 390.640 ;
        RECT 4.000 387.240 1078.020 388.640 ;
        RECT 4.000 385.240 1078.420 387.240 ;
        RECT 4.400 383.840 1078.420 385.240 ;
        RECT 4.000 378.440 1078.420 383.840 ;
        RECT 4.400 377.040 1078.020 378.440 ;
        RECT 4.000 371.640 1078.420 377.040 ;
        RECT 4.400 370.240 1078.020 371.640 ;
        RECT 4.000 364.840 1078.420 370.240 ;
        RECT 4.400 363.440 1078.020 364.840 ;
        RECT 4.000 358.040 1078.420 363.440 ;
        RECT 4.400 356.640 1078.020 358.040 ;
        RECT 4.000 351.240 1078.420 356.640 ;
        RECT 4.400 349.840 1078.020 351.240 ;
        RECT 4.000 344.440 1078.420 349.840 ;
        RECT 4.400 343.040 1078.020 344.440 ;
        RECT 4.000 337.640 1078.420 343.040 ;
        RECT 4.400 336.240 1078.020 337.640 ;
        RECT 4.000 330.840 1078.420 336.240 ;
        RECT 4.400 329.440 1078.020 330.840 ;
        RECT 4.000 324.040 1078.420 329.440 ;
        RECT 4.400 322.640 1078.020 324.040 ;
        RECT 4.000 317.240 1078.420 322.640 ;
        RECT 4.400 315.840 1078.020 317.240 ;
        RECT 4.000 310.440 1078.420 315.840 ;
        RECT 4.400 309.040 1078.020 310.440 ;
        RECT 4.000 303.640 1078.420 309.040 ;
        RECT 4.000 302.240 1078.020 303.640 ;
        RECT 4.000 300.240 1078.420 302.240 ;
        RECT 4.400 298.840 1078.420 300.240 ;
        RECT 4.000 296.840 1078.420 298.840 ;
        RECT 4.000 295.440 1078.020 296.840 ;
        RECT 4.000 293.440 1078.420 295.440 ;
        RECT 4.400 292.040 1078.420 293.440 ;
        RECT 4.000 290.040 1078.420 292.040 ;
        RECT 4.000 288.640 1078.020 290.040 ;
        RECT 4.000 286.640 1078.420 288.640 ;
        RECT 4.400 285.240 1078.420 286.640 ;
        RECT 4.000 283.240 1078.420 285.240 ;
        RECT 4.000 281.840 1078.020 283.240 ;
        RECT 4.000 279.840 1078.420 281.840 ;
        RECT 4.400 278.440 1078.420 279.840 ;
        RECT 4.000 273.040 1078.420 278.440 ;
        RECT 4.400 271.640 1078.020 273.040 ;
        RECT 4.000 266.240 1078.420 271.640 ;
        RECT 4.400 264.840 1078.020 266.240 ;
        RECT 4.000 259.440 1078.420 264.840 ;
        RECT 4.400 258.040 1078.020 259.440 ;
        RECT 4.000 252.640 1078.420 258.040 ;
        RECT 4.400 251.240 1078.020 252.640 ;
        RECT 4.000 245.840 1078.420 251.240 ;
        RECT 4.400 244.440 1078.020 245.840 ;
        RECT 4.000 239.040 1078.420 244.440 ;
        RECT 4.400 237.640 1078.020 239.040 ;
        RECT 4.000 232.240 1078.420 237.640 ;
        RECT 4.400 230.840 1078.020 232.240 ;
        RECT 4.000 225.440 1078.420 230.840 ;
        RECT 4.400 224.040 1078.020 225.440 ;
        RECT 4.000 218.640 1078.420 224.040 ;
        RECT 4.400 217.240 1078.020 218.640 ;
        RECT 4.000 211.840 1078.420 217.240 ;
        RECT 4.400 210.440 1078.020 211.840 ;
        RECT 4.000 205.040 1078.420 210.440 ;
        RECT 4.400 203.640 1078.020 205.040 ;
        RECT 4.000 198.240 1078.420 203.640 ;
        RECT 4.000 196.840 1078.020 198.240 ;
        RECT 4.000 194.840 1078.420 196.840 ;
        RECT 4.400 193.440 1078.420 194.840 ;
        RECT 4.000 191.440 1078.420 193.440 ;
        RECT 4.000 190.040 1078.020 191.440 ;
        RECT 4.000 188.040 1078.420 190.040 ;
        RECT 4.400 186.640 1078.420 188.040 ;
        RECT 4.000 184.640 1078.420 186.640 ;
        RECT 4.000 183.240 1078.020 184.640 ;
        RECT 4.000 181.240 1078.420 183.240 ;
        RECT 4.400 179.840 1078.420 181.240 ;
        RECT 4.000 174.440 1078.420 179.840 ;
        RECT 4.400 173.040 1078.020 174.440 ;
        RECT 4.000 167.640 1078.420 173.040 ;
        RECT 4.400 166.240 1078.020 167.640 ;
        RECT 4.000 160.840 1078.420 166.240 ;
        RECT 4.400 159.440 1078.020 160.840 ;
        RECT 4.000 154.040 1078.420 159.440 ;
        RECT 4.400 152.640 1078.020 154.040 ;
        RECT 4.000 147.240 1078.420 152.640 ;
        RECT 4.400 145.840 1078.020 147.240 ;
        RECT 4.000 140.440 1078.420 145.840 ;
        RECT 4.400 139.040 1078.020 140.440 ;
        RECT 4.000 133.640 1078.420 139.040 ;
        RECT 4.400 132.240 1078.020 133.640 ;
        RECT 4.000 126.840 1078.420 132.240 ;
        RECT 4.400 125.440 1078.020 126.840 ;
        RECT 4.000 120.040 1078.420 125.440 ;
        RECT 4.400 118.640 1078.020 120.040 ;
        RECT 4.000 113.240 1078.420 118.640 ;
        RECT 4.400 111.840 1078.020 113.240 ;
        RECT 4.000 106.440 1078.420 111.840 ;
        RECT 4.400 105.040 1078.020 106.440 ;
        RECT 4.000 99.640 1078.420 105.040 ;
        RECT 4.000 98.240 1078.020 99.640 ;
        RECT 4.000 96.240 1078.420 98.240 ;
        RECT 4.400 94.840 1078.420 96.240 ;
        RECT 4.000 92.840 1078.420 94.840 ;
        RECT 4.000 91.440 1078.020 92.840 ;
        RECT 4.000 89.440 1078.420 91.440 ;
        RECT 4.400 88.040 1078.420 89.440 ;
        RECT 4.000 86.040 1078.420 88.040 ;
        RECT 4.000 84.640 1078.020 86.040 ;
        RECT 4.000 82.640 1078.420 84.640 ;
        RECT 4.400 81.240 1078.420 82.640 ;
        RECT 4.000 79.240 1078.420 81.240 ;
        RECT 4.000 77.840 1078.020 79.240 ;
        RECT 4.000 75.840 1078.420 77.840 ;
        RECT 4.400 74.440 1078.420 75.840 ;
        RECT 4.000 69.040 1078.420 74.440 ;
        RECT 4.400 67.640 1078.020 69.040 ;
        RECT 4.000 62.240 1078.420 67.640 ;
        RECT 4.400 60.840 1078.020 62.240 ;
        RECT 4.000 55.440 1078.420 60.840 ;
        RECT 4.400 54.040 1078.020 55.440 ;
        RECT 4.000 48.640 1078.420 54.040 ;
        RECT 4.400 47.240 1078.020 48.640 ;
        RECT 4.000 41.840 1078.420 47.240 ;
        RECT 4.400 40.440 1078.020 41.840 ;
        RECT 4.000 35.040 1078.420 40.440 ;
        RECT 4.400 33.640 1078.020 35.040 ;
        RECT 4.000 28.240 1078.420 33.640 ;
        RECT 4.400 26.840 1078.020 28.240 ;
        RECT 4.000 21.440 1078.420 26.840 ;
        RECT 4.400 20.040 1078.020 21.440 ;
        RECT 4.000 14.640 1078.420 20.040 ;
        RECT 4.400 13.240 1078.020 14.640 ;
        RECT 4.000 10.715 1078.420 13.240 ;
      LAYER met4 ;
        RECT 10.910 12.415 24.320 1034.785 ;
        RECT 26.720 12.415 27.620 1034.785 ;
        RECT 30.020 906.780 204.320 1034.785 ;
        RECT 206.720 907.400 207.620 1034.785 ;
        RECT 210.020 907.400 384.320 1034.785 ;
        RECT 386.720 907.400 387.620 1034.785 ;
        RECT 206.720 906.780 387.620 907.400 ;
        RECT 390.020 906.780 564.320 1034.785 ;
        RECT 30.020 490.720 564.320 906.780 ;
        RECT 30.020 456.780 204.320 490.720 ;
        RECT 206.720 490.100 384.320 490.720 ;
        RECT 206.720 457.400 207.620 490.100 ;
        RECT 210.020 457.400 384.320 490.100 ;
        RECT 386.720 457.400 387.620 490.720 ;
        RECT 206.720 456.780 387.620 457.400 ;
        RECT 390.020 456.780 564.320 490.720 ;
        RECT 30.020 40.720 564.320 456.780 ;
        RECT 30.020 12.415 204.320 40.720 ;
        RECT 206.720 40.100 384.320 40.720 ;
        RECT 206.720 12.415 207.620 40.100 ;
        RECT 210.020 12.415 384.320 40.100 ;
        RECT 386.720 12.415 387.620 40.720 ;
        RECT 390.020 12.415 564.320 40.720 ;
        RECT 566.720 12.415 567.620 1034.785 ;
        RECT 570.020 12.415 744.320 1034.785 ;
        RECT 746.720 12.415 747.620 1034.785 ;
        RECT 750.020 12.415 924.320 1034.785 ;
        RECT 926.720 12.415 927.620 1034.785 ;
        RECT 930.020 12.415 1064.145 1034.785 ;
      LAYER met5 ;
        RECT 10.700 756.580 691.260 913.700 ;
        RECT 10.700 576.580 691.260 748.480 ;
        RECT 10.700 476.700 691.260 568.480 ;
        RECT 10.700 468.500 23.120 476.700 ;
        RECT 571.220 468.500 691.260 476.700 ;
        RECT 10.700 396.580 691.260 468.500 ;
        RECT 10.700 216.580 691.260 388.480 ;
        RECT 10.700 45.100 691.260 208.480 ;
  END
END soc_now_caravel_top
END LIBRARY

