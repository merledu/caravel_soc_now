##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Tue Jun  7 02:10:49 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO soc_now_caravel_top
  CLASS BLOCK ;
  SIZE 1222.220000 BY 1061.140000 ;
  FOREIGN soc_now_caravel_top 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 66.7041 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 356.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.704 LAYER met3  ;
    ANTENNAMAXAREACAR 76.345 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 393.923 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.107277 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1.920000 0.000000 2.220000 0.800000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 77.6717 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 415.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0995 LAYER met3  ;
    ANTENNAMAXAREACAR 201.914 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1030.33 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.54952 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 59.5296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 318.432 LAYER met4  ;
    ANTENNAGATEAREA 2.4465 LAYER met4  ;
    ANTENNAMAXAREACAR 226.246 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1160.48 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.679499 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 0.480000 0.600000 0.880000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 255.380000 0.000000 255.680000 0.800000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 85.640000 0.000000 85.940000 0.800000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 257.680000 0.000000 257.980000 0.800000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 252.620000 0.000000 252.920000 0.800000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.320000 0.000000 250.620000 0.800000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 248.020000 0.000000 248.320000 0.800000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 245.260000 0.000000 245.560000 0.800000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 164.300000 0.000000 164.600000 0.800000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 162.000000 0.000000 162.300000 0.800000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 159.240000 0.000000 159.540000 0.800000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.940000 0.000000 157.240000 0.800000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 154.640000 0.000000 154.940000 0.800000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 151.880000 0.000000 152.180000 0.800000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.580000 0.000000 149.880000 0.800000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.820000 0.000000 147.120000 0.800000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 144.520000 0.000000 144.820000 0.800000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 142.220000 0.000000 142.520000 0.800000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 139.920000 0.000000 140.220000 0.800000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 137.160000 0.000000 137.460000 0.800000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 134.860000 0.000000 135.160000 0.800000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 132.100000 0.000000 132.400000 0.800000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.800000 0.000000 130.100000 0.800000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 127.500000 0.000000 127.800000 0.800000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 125.200000 0.000000 125.500000 0.800000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 122.440000 0.000000 122.740000 0.800000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 120.140000 0.000000 120.440000 0.800000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.840000 0.000000 118.140000 0.800000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.080000 0.000000 115.380000 0.800000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 112.780000 0.000000 113.080000 0.800000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.020000 0.000000 110.320000 0.800000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.720000 0.000000 108.020000 0.800000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 105.420000 0.000000 105.720000 0.800000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.660000 0.000000 102.960000 0.800000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.360000 0.000000 100.660000 0.800000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 98.060000 0.000000 98.360000 0.800000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.300000 0.000000 95.600000 0.800000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 93.000000 0.000000 93.300000 0.800000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.700000 0.000000 91.000000 0.800000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 87.940000 0.000000 88.240000 0.800000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.340000 0.000000 83.640000 0.800000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.580000 0.000000 80.880000 0.800000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.280000 0.000000 78.580000 0.800000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.980000 0.000000 76.280000 0.800000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 73.220000 0.000000 73.520000 0.800000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.920000 0.000000 71.220000 0.800000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.620000 0.000000 68.920000 0.800000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.860000 0.000000 66.160000 0.800000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 63.560000 0.000000 63.860000 0.800000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.800000 0.000000 61.100000 0.800000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.500000 0.000000 58.800000 0.800000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.200000 0.000000 56.500000 0.800000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 53.440000 0.000000 53.740000 0.800000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 51.140000 0.000000 51.440000 0.800000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 48.840000 0.000000 49.140000 0.800000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.080000 0.000000 46.380000 0.800000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 43.780000 0.000000 44.080000 0.800000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.480000 0.000000 41.780000 0.800000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 38.720000 0.000000 39.020000 0.800000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.420000 0.000000 36.720000 0.800000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 34.120000 0.000000 34.420000 0.800000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.360000 0.000000 31.660000 0.800000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 29.060000 0.000000 29.360000 0.800000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.760000 0.000000 27.060000 0.800000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.000000 0.000000 24.300000 0.800000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 21.700000 0.000000 22.000000 0.800000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 19.400000 0.000000 19.700000 0.800000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.640000 0.000000 16.940000 0.800000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 14.340000 0.000000 14.640000 0.800000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 12.040000 0.000000 12.340000 0.800000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 9.280000 0.000000 9.580000 0.800000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 6.980000 0.000000 7.280000 0.800000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.837 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.61 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 4.220000 0.000000 4.520000 0.800000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.902 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1152.07 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 242.960000 0.000000 243.260000 0.800000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 240.660000 0.000000 240.960000 0.800000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 237.900000 0.000000 238.200000 0.800000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 235.600000 0.000000 235.900000 0.800000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 233.300000 0.000000 233.600000 0.800000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 230.540000 0.000000 230.840000 0.800000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 228.240000 0.000000 228.540000 0.800000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 225.940000 0.000000 226.240000 0.800000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 223.180000 0.000000 223.480000 0.800000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 220.880000 0.000000 221.180000 0.800000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 218.580000 0.000000 218.880000 0.800000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 215.820000 0.000000 216.120000 0.800000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 213.520000 0.000000 213.820000 0.800000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1152.02 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 211.220000 0.000000 211.520000 0.800000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1152.02 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 208.460000 0.000000 208.760000 0.800000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 206.160000 0.000000 206.460000 0.800000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 203.400000 0.000000 203.700000 0.800000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 201.100000 0.000000 201.400000 0.800000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 198.800000 0.000000 199.100000 0.800000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 196.040000 0.000000 196.340000 0.800000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 193.740000 0.000000 194.040000 0.800000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 191.440000 0.000000 191.740000 0.800000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 189.140000 0.000000 189.440000 0.800000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 186.380000 0.000000 186.680000 0.800000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 184.080000 0.000000 184.380000 0.800000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 181.320000 0.000000 181.620000 0.800000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 179.020000 0.000000 179.320000 0.800000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 176.720000 0.000000 177.020000 0.800000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 173.960000 0.000000 174.260000 0.800000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 171.660000 0.000000 171.960000 0.800000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 169.360000 0.000000 169.660000 0.800000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.902 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1152.07 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 166.600000 0.000000 166.900000 0.800000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 572.320000 0.000000 572.620000 0.800000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 570.020000 0.000000 570.320000 0.800000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 567.720000 0.000000 568.020000 0.800000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 564.960000 0.000000 565.260000 0.800000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 562.660000 0.000000 562.960000 0.800000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 559.900000 0.000000 560.200000 0.800000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.600000 0.000000 557.900000 0.800000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 555.300000 0.000000 555.600000 0.800000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 553.000000 0.000000 553.300000 0.800000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 550.240000 0.000000 550.540000 0.800000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 547.940000 0.000000 548.240000 0.800000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 545.640000 0.000000 545.940000 0.800000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 542.880000 0.000000 543.180000 0.800000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 540.580000 0.000000 540.880000 0.800000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 537.820000 0.000000 538.120000 0.800000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 535.520000 0.000000 535.820000 0.800000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 533.220000 0.000000 533.520000 0.800000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 530.460000 0.000000 530.760000 0.800000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 528.160000 0.000000 528.460000 0.800000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 525.860000 0.000000 526.160000 0.800000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 523.100000 0.000000 523.400000 0.800000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 520.800000 0.000000 521.100000 0.800000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 518.500000 0.000000 518.800000 0.800000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 515.740000 0.000000 516.040000 0.800000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 513.440000 0.000000 513.740000 0.800000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 511.140000 0.000000 511.440000 0.800000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 508.380000 0.000000 508.680000 0.800000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 506.080000 0.000000 506.380000 0.800000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 503.780000 0.000000 504.080000 0.800000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 501.020000 0.000000 501.320000 0.800000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 498.720000 0.000000 499.020000 0.800000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.420000 0.000000 496.720000 0.800000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 493.660000 0.000000 493.960000 0.800000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 491.360000 0.000000 491.660000 0.800000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 489.060000 0.000000 489.360000 0.800000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.300000 0.000000 486.600000 0.800000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 484.000000 0.000000 484.300000 0.800000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 481.700000 0.000000 482.000000 0.800000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 478.940000 0.000000 479.240000 0.800000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.640000 0.000000 476.940000 0.800000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 474.340000 0.000000 474.640000 0.800000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 471.580000 0.000000 471.880000 0.800000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 469.280000 0.000000 469.580000 0.800000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 466.520000 0.000000 466.820000 0.800000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 464.220000 0.000000 464.520000 0.800000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.920000 0.000000 462.220000 0.800000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 459.160000 0.000000 459.460000 0.800000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.860000 0.000000 457.160000 0.800000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 454.560000 0.000000 454.860000 0.800000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 451.800000 0.000000 452.100000 0.800000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 449.500000 0.000000 449.800000 0.800000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 447.200000 0.000000 447.500000 0.800000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.440000 0.000000 444.740000 0.800000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 442.140000 0.000000 442.440000 0.800000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 439.840000 0.000000 440.140000 0.800000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 437.080000 0.000000 437.380000 0.800000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 434.780000 0.000000 435.080000 0.800000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 432.480000 0.000000 432.780000 0.800000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 429.720000 0.000000 430.020000 0.800000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.420000 0.000000 427.720000 0.800000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 425.120000 0.000000 425.420000 0.800000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 422.360000 0.000000 422.660000 0.800000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 420.060000 0.000000 420.360000 0.800000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 417.300000 0.000000 417.600000 0.800000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 415.000000 0.000000 415.300000 0.800000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 412.700000 0.000000 413.000000 0.800000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 409.940000 0.000000 410.240000 0.800000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 407.640000 0.000000 407.940000 0.800000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 405.340000 0.000000 405.640000 0.800000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 403.040000 0.000000 403.340000 0.800000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.280000 0.000000 400.580000 0.800000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 397.980000 0.000000 398.280000 0.800000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.220000 0.000000 395.520000 0.800000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 392.920000 0.000000 393.220000 0.800000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 390.620000 0.000000 390.920000 0.800000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 387.860000 0.000000 388.160000 0.800000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 385.560000 0.000000 385.860000 0.800000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.260000 0.000000 383.560000 0.800000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 380.500000 0.000000 380.800000 0.800000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 378.200000 0.000000 378.500000 0.800000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 375.900000 0.000000 376.200000 0.800000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 373.140000 0.000000 373.440000 0.800000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.840000 0.000000 371.140000 0.800000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.540000 0.000000 368.840000 0.800000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 365.780000 0.000000 366.080000 0.800000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 363.480000 0.000000 363.780000 0.800000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 361.180000 0.000000 361.480000 0.800000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 358.420000 0.000000 358.720000 0.800000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.120000 0.000000 356.420000 0.800000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 353.820000 0.000000 354.120000 0.800000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 351.060000 0.000000 351.360000 0.800000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 348.760000 0.000000 349.060000 0.800000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000000 0.000000 346.300000 0.800000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 343.700000 0.000000 344.000000 0.800000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 341.400000 0.000000 341.700000 0.800000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 339.100000 0.000000 339.400000 0.800000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 336.340000 0.000000 336.640000 0.800000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 334.040000 0.000000 334.340000 0.800000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 331.740000 0.000000 332.040000 0.800000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 328.980000 0.000000 329.280000 0.800000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 326.680000 0.000000 326.980000 0.800000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 323.920000 0.000000 324.220000 0.800000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 321.620000 0.000000 321.920000 0.800000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 319.320000 0.000000 319.620000 0.800000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 316.560000 0.000000 316.860000 0.800000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 314.260000 0.000000 314.560000 0.800000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 311.960000 0.000000 312.260000 0.800000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 309.200000 0.000000 309.500000 0.800000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 306.900000 0.000000 307.200000 0.800000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 304.600000 0.000000 304.900000 0.800000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 301.840000 0.000000 302.140000 0.800000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 299.540000 0.000000 299.840000 0.800000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 18.9183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 77.8115 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 297.240000 0.000000 297.540000 0.800000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 18.2917 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 80.8909 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 294.480000 0.000000 294.780000 0.800000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 16.4437 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 65.621 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 292.180000 0.000000 292.480000 0.800000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 12.0035 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.5826 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.396701 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 289.880000 0.000000 290.180000 0.800000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 11.3974 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 53.6879 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 287.120000 0.000000 287.420000 0.800000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7292 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 16.6965 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 80.2313 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 284.820000 0.000000 285.120000 0.800000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 6.51939 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 31.5657 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 282.520000 0.000000 282.820000 0.800000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 6.04505 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.4646 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.24303 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 279.760000 0.000000 280.060000 0.800000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 11.0904 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 52.1004 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 277.460000 0.000000 277.760000 0.800000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 7.81455 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.9202 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 274.700000 0.000000 275.000000 0.800000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 6.42823 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 28.7896 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 272.400000 0.000000 272.700000 0.800000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 7.56848 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.6899 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.288485 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 270.100000 0.000000 270.400000 0.800000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 5.15163 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 21.8325 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.335662 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 267.340000 0.000000 267.640000 0.800000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 8.96101 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.2919 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 265.040000 0.000000 265.340000 0.800000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.80256 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 24.0317 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.261549 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 262.740000 0.000000 263.040000 0.800000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 8.29554 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.1208 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 259.980000 0.000000 260.280000 0.800000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.4005 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.1959 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 366.697 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.828 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.644 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 886.960000 0.000000 887.260000 0.800000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.0967 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 365.557 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 410.504 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 884.660000 0.000000 884.960000 0.800000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.0967 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 365.557 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 410.504 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 882.360000 0.000000 882.660000 0.800000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.0967 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 365.557 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 410.504 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 879.600000 0.000000 879.900000 0.800000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.0967 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 365.557 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 410.504 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 877.300000 0.000000 877.600000 0.800000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.0967 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 365.557 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 410.504 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 875.000000 0.000000 875.300000 0.800000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.0967 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 366.453 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.4 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 872.240000 0.000000 872.540000 0.800000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.0967 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 366.453 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.4 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 869.940000 0.000000 870.240000 0.800000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.0967 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 366.453 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.4 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 867.640000 0.000000 867.940000 0.800000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 68.0967 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 366.453 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.4 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 864.880000 0.000000 865.180000 0.800000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 78.484 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 410.31 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 85.116 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 455.257 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 862.580000 0.000000 862.880000 0.800000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.291 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 67.6387 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 360.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 74.2707 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 405.618 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 860.280000 0.000000 860.580000 0.800000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2923 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.63 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 857.520000 0.000000 857.820000 0.800000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 855.220000 0.000000 855.520000 0.800000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 852.920000 0.000000 853.220000 0.800000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 850.160000 0.000000 850.460000 0.800000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 847.860000 0.000000 848.160000 0.800000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 845.560000 0.000000 845.860000 0.800000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 842.800000 0.000000 843.100000 0.800000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 840.500000 0.000000 840.800000 0.800000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 838.200000 0.000000 838.500000 0.800000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 835.440000 0.000000 835.740000 0.800000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 833.140000 0.000000 833.440000 0.800000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 830.840000 0.000000 831.140000 0.800000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 828.080000 0.000000 828.380000 0.800000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 825.780000 0.000000 826.080000 0.800000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 823.020000 0.000000 823.320000 0.800000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 820.720000 0.000000 821.020000 0.800000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 818.420000 0.000000 818.720000 0.800000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 816.120000 0.000000 816.420000 0.800000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 813.360000 0.000000 813.660000 0.800000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 811.060000 0.000000 811.360000 0.800000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 808.300000 0.000000 808.600000 0.800000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 806.000000 0.000000 806.300000 0.800000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 803.700000 0.000000 804.000000 0.800000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 800.940000 0.000000 801.240000 0.800000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 798.640000 0.000000 798.940000 0.800000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 796.340000 0.000000 796.640000 0.800000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 793.580000 0.000000 793.880000 0.800000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 791.280000 0.000000 791.580000 0.800000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 788.980000 0.000000 789.280000 0.800000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 786.220000 0.000000 786.520000 0.800000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 783.920000 0.000000 784.220000 0.800000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 781.620000 0.000000 781.920000 0.800000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 778.860000 0.000000 779.160000 0.800000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 776.560000 0.000000 776.860000 0.800000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 773.800000 0.000000 774.100000 0.800000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 771.500000 0.000000 771.800000 0.800000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 769.200000 0.000000 769.500000 0.800000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 766.900000 0.000000 767.200000 0.800000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 764.140000 0.000000 764.440000 0.800000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 761.840000 0.000000 762.140000 0.800000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 759.540000 0.000000 759.840000 0.800000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 756.780000 0.000000 757.080000 0.800000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 754.480000 0.000000 754.780000 0.800000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 751.720000 0.000000 752.020000 0.800000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 749.420000 0.000000 749.720000 0.800000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 747.120000 0.000000 747.420000 0.800000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 744.360000 0.000000 744.660000 0.800000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 742.060000 0.000000 742.360000 0.800000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 739.760000 0.000000 740.060000 0.800000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 737.000000 0.000000 737.300000 0.800000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 734.700000 0.000000 735.000000 0.800000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 732.400000 0.000000 732.700000 0.800000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 729.640000 0.000000 729.940000 0.800000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 727.340000 0.000000 727.640000 0.800000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 725.040000 0.000000 725.340000 0.800000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 722.280000 0.000000 722.580000 0.800000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 719.980000 0.000000 720.280000 0.800000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 717.680000 0.000000 717.980000 0.800000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 714.920000 0.000000 715.220000 0.800000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 712.620000 0.000000 712.920000 0.800000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 710.320000 0.000000 710.620000 0.800000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1636.58 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 707.560000 0.000000 707.860000 0.800000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 705.260000 0.000000 705.560000 0.800000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 702.960000 0.000000 703.260000 0.800000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 700.200000 0.000000 700.500000 0.800000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 697.900000 0.000000 698.200000 0.800000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 695.600000 0.000000 695.900000 0.800000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 692.840000 0.000000 693.140000 0.800000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 690.540000 0.000000 690.840000 0.800000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 688.240000 0.000000 688.540000 0.800000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 685.480000 0.000000 685.780000 0.800000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1637.41 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 683.180000 0.000000 683.480000 0.800000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.2728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 316.795 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1683.97 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.429108 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 680.420000 0.000000 680.720000 0.800000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 65.1828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 347.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.213 LAYER met3  ;
    ANTENNAMAXAREACAR 306.023 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1632.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 678.120000 0.000000 678.420000 0.800000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.902 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1152.07 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 675.820000 0.000000 676.120000 0.800000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 673.060000 0.000000 673.360000 0.800000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 670.760000 0.000000 671.060000 0.800000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1152.02 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 668.460000 0.000000 668.760000 0.800000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1152.02 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 665.700000 0.000000 666.000000 0.800000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 663.400000 0.000000 663.700000 0.800000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 661.100000 0.000000 661.400000 0.800000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 658.340000 0.000000 658.640000 0.800000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 656.040000 0.000000 656.340000 0.800000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 653.740000 0.000000 654.040000 0.800000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 650.980000 0.000000 651.280000 0.800000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 648.680000 0.000000 648.980000 0.800000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 646.380000 0.000000 646.680000 0.800000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 643.620000 0.000000 643.920000 0.800000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 641.320000 0.000000 641.620000 0.800000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 639.020000 0.000000 639.320000 0.800000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 636.260000 0.000000 636.560000 0.800000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 633.960000 0.000000 634.260000 0.800000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 631.200000 0.000000 631.500000 0.800000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 628.900000 0.000000 629.200000 0.800000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 626.600000 0.000000 626.900000 0.800000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1152.02 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 623.840000 0.000000 624.140000 0.800000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1152.02 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 621.540000 0.000000 621.840000 0.800000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 619.240000 0.000000 619.540000 0.800000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 616.940000 0.000000 617.240000 0.800000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 614.180000 0.000000 614.480000 0.800000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 611.880000 0.000000 612.180000 0.800000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 609.120000 0.000000 609.420000 0.800000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 606.820000 0.000000 607.120000 0.800000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 604.520000 0.000000 604.820000 0.800000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 602.220000 0.000000 602.520000 0.800000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 599.460000 0.000000 599.760000 0.800000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 597.160000 0.000000 597.460000 0.800000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 594.400000 0.000000 594.700000 0.800000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 592.100000 0.000000 592.400000 0.800000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 589.800000 0.000000 590.100000 0.800000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 587.040000 0.000000 587.340000 0.800000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 584.740000 0.000000 585.040000 0.800000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 582.440000 0.000000 582.740000 0.800000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 579.680000 0.000000 579.980000 0.800000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1151.85 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 577.380000 0.000000 577.680000 0.800000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 215.792 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1150.89 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 575.080000 0.000000 575.380000 0.800000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1202.060000 0.000000 1202.360000 0.800000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1199.300000 0.000000 1199.600000 0.800000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1197.000000 0.000000 1197.300000 0.800000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1194.700000 0.000000 1195.000000 0.800000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1191.940000 0.000000 1192.240000 0.800000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1189.640000 0.000000 1189.940000 0.800000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1187.340000 0.000000 1187.640000 0.800000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1184.580000 0.000000 1184.880000 0.800000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1182.280000 0.000000 1182.580000 0.800000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1179.980000 0.000000 1180.280000 0.800000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1177.220000 0.000000 1177.520000 0.800000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1174.920000 0.000000 1175.220000 0.800000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1172.620000 0.000000 1172.920000 0.800000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1169.860000 0.000000 1170.160000 0.800000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1167.560000 0.000000 1167.860000 0.800000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1164.800000 0.000000 1165.100000 0.800000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1162.500000 0.000000 1162.800000 0.800000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1160.200000 0.000000 1160.500000 0.800000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1157.440000 0.000000 1157.740000 0.800000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1155.140000 0.000000 1155.440000 0.800000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1152.840000 0.000000 1153.140000 0.800000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1150.080000 0.000000 1150.380000 0.800000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1147.780000 0.000000 1148.080000 0.800000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1145.480000 0.000000 1145.780000 0.800000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1142.720000 0.000000 1143.020000 0.800000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1140.420000 0.000000 1140.720000 0.800000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1138.120000 0.000000 1138.420000 0.800000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1135.360000 0.000000 1135.660000 0.800000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1133.060000 0.000000 1133.360000 0.800000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1130.760000 0.000000 1131.060000 0.800000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1128.000000 0.000000 1128.300000 0.800000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1125.700000 0.000000 1126.000000 0.800000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1123.400000 0.000000 1123.700000 0.800000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1120.640000 0.000000 1120.940000 0.800000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1118.340000 0.000000 1118.640000 0.800000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1116.040000 0.000000 1116.340000 0.800000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1113.280000 0.000000 1113.580000 0.800000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1110.980000 0.000000 1111.280000 0.800000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1108.680000 0.000000 1108.980000 0.800000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1105.920000 0.000000 1106.220000 0.800000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1103.620000 0.000000 1103.920000 0.800000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1101.320000 0.000000 1101.620000 0.800000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1098.560000 0.000000 1098.860000 0.800000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.260000 0.000000 1096.560000 0.800000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1093.500000 0.000000 1093.800000 0.800000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1091.200000 0.000000 1091.500000 0.800000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1088.900000 0.000000 1089.200000 0.800000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1086.140000 0.000000 1086.440000 0.800000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1083.840000 0.000000 1084.140000 0.800000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1081.540000 0.000000 1081.840000 0.800000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1079.240000 0.000000 1079.540000 0.800000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1076.480000 0.000000 1076.780000 0.800000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1074.180000 0.000000 1074.480000 0.800000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1071.420000 0.000000 1071.720000 0.800000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1069.120000 0.000000 1069.420000 0.800000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1066.820000 0.000000 1067.120000 0.800000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1064.060000 0.000000 1064.360000 0.800000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1061.760000 0.000000 1062.060000 0.800000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1059.460000 0.000000 1059.760000 0.800000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1056.700000 0.000000 1057.000000 0.800000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1054.400000 0.000000 1054.700000 0.800000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1052.100000 0.000000 1052.400000 0.800000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1049.340000 0.000000 1049.640000 0.800000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1047.040000 0.000000 1047.340000 0.800000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1044.740000 0.000000 1045.040000 0.800000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1041.980000 0.000000 1042.280000 0.800000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1039.680000 0.000000 1039.980000 0.800000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1036.920000 0.000000 1037.220000 0.800000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1034.620000 0.000000 1034.920000 0.800000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1032.320000 0.000000 1032.620000 0.800000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1030.020000 0.000000 1030.320000 0.800000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1027.260000 0.000000 1027.560000 0.800000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1024.960000 0.000000 1025.260000 0.800000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1022.200000 0.000000 1022.500000 0.800000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.900000 0.000000 1020.200000 0.800000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1017.600000 0.000000 1017.900000 0.800000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1014.840000 0.000000 1015.140000 0.800000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1012.540000 0.000000 1012.840000 0.800000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1010.240000 0.000000 1010.540000 0.800000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1007.480000 0.000000 1007.780000 0.800000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1005.180000 0.000000 1005.480000 0.800000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1002.880000 0.000000 1003.180000 0.800000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1000.120000 0.000000 1000.420000 0.800000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 997.820000 0.000000 998.120000 0.800000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 995.520000 0.000000 995.820000 0.800000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 992.760000 0.000000 993.060000 0.800000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 990.460000 0.000000 990.760000 0.800000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 987.700000 0.000000 988.000000 0.800000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 985.400000 0.000000 985.700000 0.800000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 983.100000 0.000000 983.400000 0.800000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 980.800000 0.000000 981.100000 0.800000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 978.040000 0.000000 978.340000 0.800000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 975.740000 0.000000 976.040000 0.800000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 973.440000 0.000000 973.740000 0.800000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 970.680000 0.000000 970.980000 0.800000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 968.380000 0.000000 968.680000 0.800000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 966.080000 0.000000 966.380000 0.800000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 963.320000 0.000000 963.620000 0.800000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 961.020000 0.000000 961.320000 0.800000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 958.720000 0.000000 959.020000 0.800000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 955.960000 0.000000 956.260000 0.800000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 953.660000 0.000000 953.960000 0.800000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 950.900000 0.000000 951.200000 0.800000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 948.600000 0.000000 948.900000 0.800000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 946.300000 0.000000 946.600000 0.800000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 943.540000 0.000000 943.840000 0.800000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 941.240000 0.000000 941.540000 0.800000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 938.940000 0.000000 939.240000 0.800000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 936.180000 0.000000 936.480000 0.800000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.880000 0.000000 934.180000 0.800000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 931.580000 0.000000 931.880000 0.800000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 928.820000 0.000000 929.120000 0.800000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 926.520000 0.000000 926.820000 0.800000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 924.220000 0.000000 924.520000 0.800000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 921.460000 0.000000 921.760000 0.800000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 919.160000 0.000000 919.460000 0.800000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 916.860000 0.000000 917.160000 0.800000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 914.100000 0.000000 914.400000 0.800000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 911.800000 0.000000 912.100000 0.800000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 909.500000 0.000000 909.800000 0.800000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 906.740000 0.000000 907.040000 0.800000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 904.440000 0.000000 904.740000 0.800000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 902.140000 0.000000 902.440000 0.800000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 899.380000 0.000000 899.680000 0.800000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 897.080000 0.000000 897.380000 0.800000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.320000 0.000000 894.620000 0.800000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 892.020000 0.000000 892.320000 0.800000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 889.720000 0.000000 890.020000 0.800000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.88 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 67.7598 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 336.277 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.643488 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 39.520000 0.600000 39.920000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 128.294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 684.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 30.2642 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 143.841 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 98.690000 0.600000 99.090000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 138.827 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 740.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 21.1892 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 102.078 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 157.860000 0.600000 158.260000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 135.053 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 720.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 25.1625 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.282 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 236.550000 0.600000 236.950000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 145.521 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 776.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 5.7388 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 26.6485 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.403566 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 315.850000 0.600000 316.250000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 148.14 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 790.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 22.9673 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 116.73 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.782377 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 394.540000 0.600000 394.940000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 134.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 718.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9392 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 52.2997 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 271.294 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 473.840000 0.600000 474.240000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.6214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.976 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 96.5863 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 486.287 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.643488 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 552.530000 0.600000 552.930000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 107.436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 573.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 60.5524 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 312.097 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 631.830000 0.600000 632.230000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 81.8836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 436.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 99.4008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 530.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 239.172 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1257.12 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 710.520000 0.600000 710.920000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.9744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 346.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 87.4628 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 442.913 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 789.210000 0.600000 789.610000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3901 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.576 LAYER met3  ;
    ANTENNAMAXAREACAR 23.9574 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 119.979 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.515823 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 31.6864 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 161.871 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 868.510000 0.600000 868.910000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 108.008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 576.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 168.878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 901.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 284.985 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1508.75 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 947.200000 0.600000 947.600000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 114.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 611.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 200.258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1068.51 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 353.713 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1803 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.782377 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1025.890000 0.600000 1026.290000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 95.6344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 510.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.5986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 40.8938 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 213.314 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 69.080000 1060.340000 69.380000 1061.140000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.8334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 109.196 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 582.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 213.424 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1082.88 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 208.000000 1060.340000 208.300000 1061.140000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 114.845 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 612.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 210.212 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1047.45 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.782377 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 346.460000 1060.340000 346.760000 1061.140000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 237.089 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1264.94 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 357.275 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1864.47 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 484.920000 1060.340000 485.220000 1061.140000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.7492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 124.13 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 662.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 223.642 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1181.56 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 623.380000 1060.340000 623.680000 1061.140000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 122.372 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 653.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 192.245 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1003.2 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 761.840000 1060.340000 762.140000 1061.140000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 121.568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 648.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 186.266 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 949.663 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.375376 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 900.300000 1060.340000 900.600000 1061.140000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.7574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 128.498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 685.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 196.042 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1031.84 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1038.760000 1060.340000 1039.060000 1061.140000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.5894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 133.757 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 713.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 222.113 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1107.59 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1177.680000 1060.340000 1177.980000 1061.140000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 194.879 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1039.34 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 213.179 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1137.42 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 330.499 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1689.91 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.782377 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 1005.150000 1222.220000 1005.550000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 119.165 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 636.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 194.323 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1023.29 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700468 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 924.630000 1222.220000 925.030000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 63.2284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 337.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 537.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 158.198 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 819.924 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 844.110000 1222.220000 844.510000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.9974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.0208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 331.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 106.862 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 555.961 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.751262 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 763.590000 1222.220000 763.990000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 190.323 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1015.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 70.2078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 374.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 113.738 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 600.485 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521897 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 683.070000 1222.220000 683.470000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4454 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.5454 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 75.3783 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 376.386 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.960948 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 603.160000 1222.220000 603.560000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 71.8788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 383.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 121.306 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 596.49 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536379 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 522.640000 1222.220000 523.040000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.7518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met4  ;
    ANTENNAMAXAREACAR 69.6461 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 348.434 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.929833 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 442.120000 1222.220000 442.520000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.702 LAYER met3  ;
    ANTENNAMAXAREACAR 79.1248 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 386.763 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.464917 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 361.600000 1222.220000 362.000000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.6403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 179.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.6134 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 43.1612 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 228.356 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854141 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 301.210000 1222.220000 301.610000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 240.820000 1222.220000 241.220000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 180.430000 1222.220000 180.830000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 120.040000 1222.220000 120.440000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 59.650000 1222.220000 60.050000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.790000 0.000000 1222.190000 0.600000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 101.744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 542.632 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 20.000000 0.600000 20.400000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 133.985 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 714.584 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 79.170000 0.600000 79.570000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 99.6714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 531.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 138.340000 0.600000 138.740000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 217.030000 0.600000 217.430000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 122.528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 653.48 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 296.330000 0.600000 296.730000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 119.023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 635.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 375.020000 0.600000 375.420000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 72.2382 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 385.736 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 453.710000 0.600000 454.110000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 139.299 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 743.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.6614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 36.8937 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 198.105 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 533.010000 0.600000 533.410000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.8088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 133.286 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 702.976 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 611.700000 0.600000 612.100000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 124.13 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 662.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 71.5206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 382.384 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 691.000000 0.600000 691.400000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 75.2656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 401.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 127.583 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 680.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 769.690000 0.600000 770.090000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 107.132 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 571.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 158.36 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 845.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 220.416 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1168.03 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.409697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 848.380000 0.600000 848.780000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 89.7676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 478.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 165.656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 883.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 250.332 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1326.52 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.571313 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 927.680000 0.600000 928.080000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 83.5576 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 445.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 196.964 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1050.94 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 274.402 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1459.28 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.409697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1006.370000 0.600000 1006.770000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 82.0974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 437.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 34.580000 1060.340000 34.880000 1061.140000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 139.23 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 744.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 162.334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 860.085 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 173.040000 1060.340000 173.340000 1061.140000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 133.169 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 710.704 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 311.960000 1060.340000 312.260000 1061.140000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 121.745 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 649.776 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 450.420000 1060.340000 450.720000 1061.140000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 103.427 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 552.08 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 588.880000 1060.340000 589.180000 1061.140000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 57.5356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 306.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 163.22 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 870.976 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 727.340000 1060.340000 727.640000 1061.140000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.2584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 177.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 118.895 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 634.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 169.167 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 898.707 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 865.800000 1060.340000 866.100000 1061.140000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1942 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 121.004 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 645.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 180.626 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 957.215 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1004.260000 1060.340000 1004.560000 1061.140000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 115.322 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 615.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 175.651 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 931.073 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.40633 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1142.720000 1060.340000 1143.020000 1061.140000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 203.939 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1087.66 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 205.804 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1098.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 290.179 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1543.51 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.40633 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 1025.280000 1222.220000 1025.680000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.8478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 484.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 134.489 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 711.941 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 944.760000 1222.220000 945.160000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.6374 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 66.7285 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 352.967 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692525 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 864.240000 1222.220000 864.640000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 72.3094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 386.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.6418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 318.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 131.001 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 684.56 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.315421 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 783.720000 1222.220000 784.120000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 85.3792 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 456.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.9708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 341.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 127.386 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 667.972 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.67569 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 703.200000 1222.220000 703.600000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 622.680000 1222.220000 623.080000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.6264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 281.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.6268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 104.075 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 545.988 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.40633 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 542.770000 1222.220000 543.170000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 54.9004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 293.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.6288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 339.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 278.958 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1483.46 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 462.250000 1222.220000 462.650000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.5948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.976 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 381.730000 1222.220000 382.130000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 321.340000 1222.220000 321.740000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9522 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 260.950000 1222.220000 261.350000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9822 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 200.560000 1222.220000 200.960000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 140.170000 1222.220000 140.570000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 79.780000 1222.220000 80.180000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 19.390000 1222.220000 19.790000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1.000000 0.000000 1.300000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 97.4214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 519.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.040000 0.600000 59.440000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 118.210000 0.600000 118.610000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 197.510000 0.600000 197.910000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 139.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 743.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 276.200000 0.600000 276.600000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 137.602 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 734.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 355.500000 0.600000 355.900000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 73.5252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 392.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 434.190000 0.600000 434.590000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 116.671 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 622.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 512.880000 0.600000 513.280000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.0434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.56 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 592.180000 0.600000 592.580000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.4804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 670.870000 0.600000 671.270000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.1114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 750.170000 0.600000 750.570000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 110.531 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 589.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 828.860000 0.600000 829.260000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 111.59 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 595.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 907.550000 0.600000 907.950000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 986.850000 0.600000 987.250000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.1904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1.460000 1060.340000 1.760000 1061.140000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 138.540000 1060.340000 138.840000 1061.140000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 45.1212 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 241.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 277.000000 1060.340000 277.300000 1061.140000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.416 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 415.460000 1060.340000 415.760000 1061.140000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 554.380000 1060.340000 554.680000 1061.140000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.55935 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.2578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 412.512 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 692.840000 1060.340000 693.140000 1061.140000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5413 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.6626 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 94.2288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 503.024 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 831.300000 1060.340000 831.600000 1061.140000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.3008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 487.408 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 969.760000 1060.340000 970.060000 1061.140000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.2584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1108.220000 1060.340000 1108.520000 1061.140000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.14935 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.6438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 339.904 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 1044.800000 1222.220000 1045.200000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.4648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 413.616 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 964.890000 1222.220000 965.290000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 118.568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 632.832 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 884.370000 1222.220000 884.770000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 194.43 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1037.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.5548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.096 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 803.850000 1222.220000 804.250000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 92.053 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 491.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.3538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.024 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 723.330000 1222.220000 723.730000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.9058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.968 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 642.810000 1222.220000 643.210000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 187.259 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 998.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.6626 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.7848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.656 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 562.290000 1222.220000 562.690000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.1744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 203.592 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 482.380000 1222.220000 482.780000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 401.860000 1222.220000 402.260000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 341.470000 1222.220000 341.870000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 281.080000 1222.220000 281.480000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 220.690000 1222.220000 221.090000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 160.300000 1222.220000 160.700000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 99.910000 1222.220000 100.310000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 39.520000 1222.220000 39.920000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 177.380000 0.600000 177.780000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 256.680000 0.600000 257.080000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 335.370000 0.600000 335.770000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 414.670000 0.600000 415.070000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 493.360000 0.600000 493.760000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 572.050000 0.600000 572.450000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 651.350000 0.600000 651.750000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 730.040000 0.600000 730.440000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 809.340000 0.600000 809.740000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 888.030000 0.600000 888.430000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 966.720000 0.600000 967.120000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1045.410000 0.600000 1045.810000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 104.040000 1060.340000 104.340000 1061.140000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 242.500000 1060.340000 242.800000 1061.140000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 380.960000 1060.340000 381.260000 1061.140000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 519.420000 1060.340000 519.720000 1061.140000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 657.880000 1060.340000 658.180000 1061.140000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.800000 1060.340000 797.100000 1061.140000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 935.260000 1060.340000 935.560000 1061.140000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1073.720000 1060.340000 1074.020000 1061.140000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1211.260000 1060.340000 1211.560000 1061.140000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 985.020000 1222.220000 985.420000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 904.500000 1222.220000 904.900000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 823.980000 1222.220000 824.380000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 743.460000 1222.220000 743.860000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 662.940000 1222.220000 663.340000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 583.030000 1222.220000 583.430000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 502.510000 1222.220000 502.910000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.620000 421.990000 1222.220000 422.390000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1204.360000 0.000000 1204.660000 0.800000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9822 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1209.420000 0.000000 1209.720000 0.800000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9372 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1211.260000 0.000000 1211.560000 0.800000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.8922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 6.63206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9466 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1206.660000 0.000000 1206.960000 0.800000 ;
    END
  END user_irq[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 7.840000 7.680000 1214.380000 9.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.840000 1051.520000 1214.380000 1053.120000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1212.780000 7.680000 1214.380000 1053.120000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.840000 7.680000 9.440000 1053.120000 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.640000 4.480000 6.240000 1056.320000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 607.250000 143.290000 608.990000 531.270000 ;
      LAYER met4 ;
        RECT 1075.770000 143.290000 1077.510000 531.270000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 607.250000 591.790000 608.990000 979.770000 ;
      LAYER met4 ;
        RECT 1075.770000 591.790000 1077.510000 979.770000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 4.640000 4.480000 1217.580000 6.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.640000 1054.720000 1217.580000 1056.320000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1215.980000 4.480000 1217.580000 1056.320000 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.640000 4.480000 6.240000 1056.320000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1079.170000 139.890000 1080.910000 534.670000 ;
      LAYER met4 ;
        RECT 603.850000 139.890000 605.590000 534.670000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'


# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 1079.170000 588.390000 1080.910000 983.170000 ;
      LAYER met4 ;
        RECT 603.850000 588.390000 605.590000 983.170000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1222.220000 1061.140000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1222.220000 1061.140000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 1222.220000 1061.140000 ;
    LAYER met3 ;
      RECT 1211.860000 1060.040000 1222.220000 1061.140000 ;
      RECT 1178.280000 1060.040000 1210.960000 1061.140000 ;
      RECT 1143.320000 1060.040000 1177.380000 1061.140000 ;
      RECT 1108.820000 1060.040000 1142.420000 1061.140000 ;
      RECT 1074.320000 1060.040000 1107.920000 1061.140000 ;
      RECT 1039.360000 1060.040000 1073.420000 1061.140000 ;
      RECT 1004.860000 1060.040000 1038.460000 1061.140000 ;
      RECT 970.360000 1060.040000 1003.960000 1061.140000 ;
      RECT 935.860000 1060.040000 969.460000 1061.140000 ;
      RECT 900.900000 1060.040000 934.960000 1061.140000 ;
      RECT 866.400000 1060.040000 900.000000 1061.140000 ;
      RECT 831.900000 1060.040000 865.500000 1061.140000 ;
      RECT 797.400000 1060.040000 831.000000 1061.140000 ;
      RECT 762.440000 1060.040000 796.500000 1061.140000 ;
      RECT 727.940000 1060.040000 761.540000 1061.140000 ;
      RECT 693.440000 1060.040000 727.040000 1061.140000 ;
      RECT 658.480000 1060.040000 692.540000 1061.140000 ;
      RECT 623.980000 1060.040000 657.580000 1061.140000 ;
      RECT 589.480000 1060.040000 623.080000 1061.140000 ;
      RECT 554.980000 1060.040000 588.580000 1061.140000 ;
      RECT 520.020000 1060.040000 554.080000 1061.140000 ;
      RECT 485.520000 1060.040000 519.120000 1061.140000 ;
      RECT 451.020000 1060.040000 484.620000 1061.140000 ;
      RECT 416.060000 1060.040000 450.120000 1061.140000 ;
      RECT 381.560000 1060.040000 415.160000 1061.140000 ;
      RECT 347.060000 1060.040000 380.660000 1061.140000 ;
      RECT 312.560000 1060.040000 346.160000 1061.140000 ;
      RECT 277.600000 1060.040000 311.660000 1061.140000 ;
      RECT 243.100000 1060.040000 276.700000 1061.140000 ;
      RECT 208.600000 1060.040000 242.200000 1061.140000 ;
      RECT 173.640000 1060.040000 207.700000 1061.140000 ;
      RECT 139.140000 1060.040000 172.740000 1061.140000 ;
      RECT 104.640000 1060.040000 138.240000 1061.140000 ;
      RECT 69.680000 1060.040000 103.740000 1061.140000 ;
      RECT 35.180000 1060.040000 68.780000 1061.140000 ;
      RECT 2.060000 1060.040000 34.280000 1061.140000 ;
      RECT 0.000000 1060.040000 1.160000 1061.140000 ;
      RECT 0.000000 1056.620000 1222.220000 1060.040000 ;
      RECT 1217.880000 1054.420000 1222.220000 1056.620000 ;
      RECT 0.000000 1054.420000 4.340000 1056.620000 ;
      RECT 0.000000 1053.420000 1222.220000 1054.420000 ;
      RECT 1214.680000 1051.220000 1222.220000 1053.420000 ;
      RECT 0.000000 1051.220000 7.540000 1053.420000 ;
      RECT 0.000000 1046.110000 1222.220000 1051.220000 ;
      RECT 0.900000 1045.500000 1222.220000 1046.110000 ;
      RECT 0.900000 1045.110000 1221.320000 1045.500000 ;
      RECT 0.000000 1044.500000 1221.320000 1045.110000 ;
      RECT 0.000000 1026.590000 1222.220000 1044.500000 ;
      RECT 0.900000 1025.980000 1222.220000 1026.590000 ;
      RECT 0.900000 1025.590000 1221.320000 1025.980000 ;
      RECT 0.000000 1024.980000 1221.320000 1025.590000 ;
      RECT 0.000000 1007.070000 1222.220000 1024.980000 ;
      RECT 0.900000 1006.070000 1222.220000 1007.070000 ;
      RECT 0.000000 1005.850000 1222.220000 1006.070000 ;
      RECT 0.000000 1004.850000 1221.320000 1005.850000 ;
      RECT 0.000000 987.550000 1222.220000 1004.850000 ;
      RECT 0.900000 986.550000 1222.220000 987.550000 ;
      RECT 0.000000 985.720000 1222.220000 986.550000 ;
      RECT 0.000000 984.720000 1221.320000 985.720000 ;
      RECT 0.000000 967.420000 1222.220000 984.720000 ;
      RECT 0.900000 966.420000 1222.220000 967.420000 ;
      RECT 0.000000 965.590000 1222.220000 966.420000 ;
      RECT 0.000000 964.590000 1221.320000 965.590000 ;
      RECT 0.000000 947.900000 1222.220000 964.590000 ;
      RECT 0.900000 946.900000 1222.220000 947.900000 ;
      RECT 0.000000 945.460000 1222.220000 946.900000 ;
      RECT 0.000000 944.460000 1221.320000 945.460000 ;
      RECT 0.000000 928.380000 1222.220000 944.460000 ;
      RECT 0.900000 927.380000 1222.220000 928.380000 ;
      RECT 0.000000 925.330000 1222.220000 927.380000 ;
      RECT 0.000000 924.330000 1221.320000 925.330000 ;
      RECT 0.000000 908.250000 1222.220000 924.330000 ;
      RECT 0.900000 907.250000 1222.220000 908.250000 ;
      RECT 0.000000 905.200000 1222.220000 907.250000 ;
      RECT 0.000000 904.200000 1221.320000 905.200000 ;
      RECT 0.000000 888.730000 1222.220000 904.200000 ;
      RECT 0.900000 887.730000 1222.220000 888.730000 ;
      RECT 0.000000 885.070000 1222.220000 887.730000 ;
      RECT 0.000000 884.070000 1221.320000 885.070000 ;
      RECT 0.000000 869.210000 1222.220000 884.070000 ;
      RECT 0.900000 868.210000 1222.220000 869.210000 ;
      RECT 0.000000 864.940000 1222.220000 868.210000 ;
      RECT 0.000000 863.940000 1221.320000 864.940000 ;
      RECT 0.000000 849.080000 1222.220000 863.940000 ;
      RECT 0.900000 848.080000 1222.220000 849.080000 ;
      RECT 0.000000 844.810000 1222.220000 848.080000 ;
      RECT 0.000000 843.810000 1221.320000 844.810000 ;
      RECT 0.000000 829.560000 1222.220000 843.810000 ;
      RECT 0.900000 828.560000 1222.220000 829.560000 ;
      RECT 0.000000 824.680000 1222.220000 828.560000 ;
      RECT 0.000000 823.680000 1221.320000 824.680000 ;
      RECT 0.000000 810.040000 1222.220000 823.680000 ;
      RECT 0.900000 809.040000 1222.220000 810.040000 ;
      RECT 0.000000 804.550000 1222.220000 809.040000 ;
      RECT 0.000000 803.550000 1221.320000 804.550000 ;
      RECT 0.000000 789.910000 1222.220000 803.550000 ;
      RECT 0.900000 788.910000 1222.220000 789.910000 ;
      RECT 0.000000 784.420000 1222.220000 788.910000 ;
      RECT 0.000000 783.420000 1221.320000 784.420000 ;
      RECT 0.000000 770.390000 1222.220000 783.420000 ;
      RECT 0.900000 769.390000 1222.220000 770.390000 ;
      RECT 0.000000 764.290000 1222.220000 769.390000 ;
      RECT 0.000000 763.290000 1221.320000 764.290000 ;
      RECT 0.000000 750.870000 1222.220000 763.290000 ;
      RECT 0.900000 749.870000 1222.220000 750.870000 ;
      RECT 0.000000 744.160000 1222.220000 749.870000 ;
      RECT 0.000000 743.160000 1221.320000 744.160000 ;
      RECT 0.000000 730.740000 1222.220000 743.160000 ;
      RECT 0.900000 729.740000 1222.220000 730.740000 ;
      RECT 0.000000 724.030000 1222.220000 729.740000 ;
      RECT 0.000000 723.030000 1221.320000 724.030000 ;
      RECT 0.000000 711.220000 1222.220000 723.030000 ;
      RECT 0.900000 710.220000 1222.220000 711.220000 ;
      RECT 0.000000 703.900000 1222.220000 710.220000 ;
      RECT 0.000000 702.900000 1221.320000 703.900000 ;
      RECT 0.000000 691.700000 1222.220000 702.900000 ;
      RECT 0.900000 690.700000 1222.220000 691.700000 ;
      RECT 0.000000 683.770000 1222.220000 690.700000 ;
      RECT 0.000000 682.770000 1221.320000 683.770000 ;
      RECT 0.000000 671.570000 1222.220000 682.770000 ;
      RECT 0.900000 670.570000 1222.220000 671.570000 ;
      RECT 0.000000 663.640000 1222.220000 670.570000 ;
      RECT 0.000000 662.640000 1221.320000 663.640000 ;
      RECT 0.000000 652.050000 1222.220000 662.640000 ;
      RECT 0.900000 651.050000 1222.220000 652.050000 ;
      RECT 0.000000 643.510000 1222.220000 651.050000 ;
      RECT 0.000000 642.510000 1221.320000 643.510000 ;
      RECT 0.000000 632.530000 1222.220000 642.510000 ;
      RECT 0.900000 631.530000 1222.220000 632.530000 ;
      RECT 0.000000 623.380000 1222.220000 631.530000 ;
      RECT 0.000000 622.380000 1221.320000 623.380000 ;
      RECT 0.000000 612.400000 1222.220000 622.380000 ;
      RECT 0.900000 611.400000 1222.220000 612.400000 ;
      RECT 0.000000 603.860000 1222.220000 611.400000 ;
      RECT 0.000000 602.860000 1221.320000 603.860000 ;
      RECT 0.000000 592.880000 1222.220000 602.860000 ;
      RECT 0.900000 591.880000 1222.220000 592.880000 ;
      RECT 0.000000 583.730000 1222.220000 591.880000 ;
      RECT 0.000000 582.730000 1221.320000 583.730000 ;
      RECT 0.000000 572.750000 1222.220000 582.730000 ;
      RECT 0.900000 571.750000 1222.220000 572.750000 ;
      RECT 0.000000 562.990000 1222.220000 571.750000 ;
      RECT 0.000000 561.990000 1221.320000 562.990000 ;
      RECT 0.000000 553.230000 1222.220000 561.990000 ;
      RECT 0.900000 552.230000 1222.220000 553.230000 ;
      RECT 0.000000 543.470000 1222.220000 552.230000 ;
      RECT 0.000000 542.470000 1221.320000 543.470000 ;
      RECT 0.000000 533.710000 1222.220000 542.470000 ;
      RECT 0.900000 532.710000 1222.220000 533.710000 ;
      RECT 0.000000 523.340000 1222.220000 532.710000 ;
      RECT 0.000000 522.340000 1221.320000 523.340000 ;
      RECT 0.000000 513.580000 1222.220000 522.340000 ;
      RECT 0.900000 512.580000 1222.220000 513.580000 ;
      RECT 0.000000 503.210000 1222.220000 512.580000 ;
      RECT 0.000000 502.210000 1221.320000 503.210000 ;
      RECT 0.000000 494.060000 1222.220000 502.210000 ;
      RECT 0.900000 493.060000 1222.220000 494.060000 ;
      RECT 0.000000 483.080000 1222.220000 493.060000 ;
      RECT 0.000000 482.080000 1221.320000 483.080000 ;
      RECT 0.000000 474.540000 1222.220000 482.080000 ;
      RECT 0.900000 473.540000 1222.220000 474.540000 ;
      RECT 0.000000 462.950000 1222.220000 473.540000 ;
      RECT 0.000000 461.950000 1221.320000 462.950000 ;
      RECT 0.000000 454.410000 1222.220000 461.950000 ;
      RECT 0.900000 453.410000 1222.220000 454.410000 ;
      RECT 0.000000 442.820000 1222.220000 453.410000 ;
      RECT 0.000000 441.820000 1221.320000 442.820000 ;
      RECT 0.000000 434.890000 1222.220000 441.820000 ;
      RECT 0.900000 433.890000 1222.220000 434.890000 ;
      RECT 0.000000 422.690000 1222.220000 433.890000 ;
      RECT 0.000000 421.690000 1221.320000 422.690000 ;
      RECT 0.000000 415.370000 1222.220000 421.690000 ;
      RECT 0.900000 414.370000 1222.220000 415.370000 ;
      RECT 0.000000 402.560000 1222.220000 414.370000 ;
      RECT 0.000000 401.560000 1221.320000 402.560000 ;
      RECT 0.000000 395.240000 1222.220000 401.560000 ;
      RECT 0.900000 394.240000 1222.220000 395.240000 ;
      RECT 0.000000 382.430000 1222.220000 394.240000 ;
      RECT 0.000000 381.430000 1221.320000 382.430000 ;
      RECT 0.000000 375.720000 1222.220000 381.430000 ;
      RECT 0.900000 374.720000 1222.220000 375.720000 ;
      RECT 0.000000 362.300000 1222.220000 374.720000 ;
      RECT 0.000000 361.300000 1221.320000 362.300000 ;
      RECT 0.000000 356.200000 1222.220000 361.300000 ;
      RECT 0.900000 355.200000 1222.220000 356.200000 ;
      RECT 0.000000 342.170000 1222.220000 355.200000 ;
      RECT 0.000000 341.170000 1221.320000 342.170000 ;
      RECT 0.000000 336.070000 1222.220000 341.170000 ;
      RECT 0.900000 335.070000 1222.220000 336.070000 ;
      RECT 0.000000 322.040000 1222.220000 335.070000 ;
      RECT 0.000000 321.040000 1221.320000 322.040000 ;
      RECT 0.000000 316.550000 1222.220000 321.040000 ;
      RECT 0.900000 315.550000 1222.220000 316.550000 ;
      RECT 0.000000 301.910000 1222.220000 315.550000 ;
      RECT 0.000000 300.910000 1221.320000 301.910000 ;
      RECT 0.000000 297.030000 1222.220000 300.910000 ;
      RECT 0.900000 296.030000 1222.220000 297.030000 ;
      RECT 0.000000 281.780000 1222.220000 296.030000 ;
      RECT 0.000000 280.780000 1221.320000 281.780000 ;
      RECT 0.000000 276.900000 1222.220000 280.780000 ;
      RECT 0.900000 275.900000 1222.220000 276.900000 ;
      RECT 0.000000 261.650000 1222.220000 275.900000 ;
      RECT 0.000000 260.650000 1221.320000 261.650000 ;
      RECT 0.000000 257.380000 1222.220000 260.650000 ;
      RECT 0.900000 256.380000 1222.220000 257.380000 ;
      RECT 0.000000 241.520000 1222.220000 256.380000 ;
      RECT 0.000000 240.520000 1221.320000 241.520000 ;
      RECT 0.000000 237.250000 1222.220000 240.520000 ;
      RECT 0.900000 236.250000 1222.220000 237.250000 ;
      RECT 0.000000 221.390000 1222.220000 236.250000 ;
      RECT 0.000000 220.390000 1221.320000 221.390000 ;
      RECT 0.000000 217.730000 1222.220000 220.390000 ;
      RECT 0.900000 216.730000 1222.220000 217.730000 ;
      RECT 0.000000 201.260000 1222.220000 216.730000 ;
      RECT 0.000000 200.260000 1221.320000 201.260000 ;
      RECT 0.000000 198.210000 1222.220000 200.260000 ;
      RECT 0.900000 197.210000 1222.220000 198.210000 ;
      RECT 0.000000 181.130000 1222.220000 197.210000 ;
      RECT 0.000000 180.130000 1221.320000 181.130000 ;
      RECT 0.000000 178.080000 1222.220000 180.130000 ;
      RECT 0.900000 177.080000 1222.220000 178.080000 ;
      RECT 0.000000 161.000000 1222.220000 177.080000 ;
      RECT 0.000000 160.000000 1221.320000 161.000000 ;
      RECT 0.000000 158.560000 1222.220000 160.000000 ;
      RECT 0.900000 157.560000 1222.220000 158.560000 ;
      RECT 0.000000 140.870000 1222.220000 157.560000 ;
      RECT 0.000000 139.870000 1221.320000 140.870000 ;
      RECT 0.000000 139.040000 1222.220000 139.870000 ;
      RECT 0.900000 138.040000 1222.220000 139.040000 ;
      RECT 0.000000 120.740000 1222.220000 138.040000 ;
      RECT 0.000000 119.740000 1221.320000 120.740000 ;
      RECT 0.000000 118.910000 1222.220000 119.740000 ;
      RECT 0.900000 117.910000 1222.220000 118.910000 ;
      RECT 0.000000 100.610000 1222.220000 117.910000 ;
      RECT 0.000000 99.610000 1221.320000 100.610000 ;
      RECT 0.000000 99.390000 1222.220000 99.610000 ;
      RECT 0.900000 98.390000 1222.220000 99.390000 ;
      RECT 0.000000 80.480000 1222.220000 98.390000 ;
      RECT 0.000000 79.870000 1221.320000 80.480000 ;
      RECT 0.900000 79.480000 1221.320000 79.870000 ;
      RECT 0.900000 78.870000 1222.220000 79.480000 ;
      RECT 0.000000 60.350000 1222.220000 78.870000 ;
      RECT 0.000000 59.740000 1221.320000 60.350000 ;
      RECT 0.900000 59.350000 1221.320000 59.740000 ;
      RECT 0.900000 58.740000 1222.220000 59.350000 ;
      RECT 0.000000 40.220000 1222.220000 58.740000 ;
      RECT 0.900000 39.220000 1221.320000 40.220000 ;
      RECT 0.000000 20.700000 1222.220000 39.220000 ;
      RECT 0.900000 20.090000 1222.220000 20.700000 ;
      RECT 0.900000 19.700000 1221.320000 20.090000 ;
      RECT 0.000000 19.090000 1221.320000 19.700000 ;
      RECT 0.000000 9.580000 1222.220000 19.090000 ;
      RECT 1214.680000 7.380000 1222.220000 9.580000 ;
      RECT 0.000000 7.380000 7.540000 9.580000 ;
      RECT 0.000000 6.380000 1222.220000 7.380000 ;
      RECT 1217.880000 4.180000 1222.220000 6.380000 ;
      RECT 0.000000 4.180000 4.340000 6.380000 ;
      RECT 0.000000 1.180000 1222.220000 4.180000 ;
      RECT 0.900000 1.100000 1222.220000 1.180000 ;
      RECT 1211.860000 0.900000 1222.220000 1.100000 ;
      RECT 1211.860000 0.000000 1221.490000 0.900000 ;
      RECT 1210.020000 0.000000 1210.960000 1.100000 ;
      RECT 1207.260000 0.000000 1209.120000 1.100000 ;
      RECT 1204.960000 0.000000 1206.360000 1.100000 ;
      RECT 1202.660000 0.000000 1204.060000 1.100000 ;
      RECT 1199.900000 0.000000 1201.760000 1.100000 ;
      RECT 1197.600000 0.000000 1199.000000 1.100000 ;
      RECT 1195.300000 0.000000 1196.700000 1.100000 ;
      RECT 1192.540000 0.000000 1194.400000 1.100000 ;
      RECT 1190.240000 0.000000 1191.640000 1.100000 ;
      RECT 1187.940000 0.000000 1189.340000 1.100000 ;
      RECT 1185.180000 0.000000 1187.040000 1.100000 ;
      RECT 1182.880000 0.000000 1184.280000 1.100000 ;
      RECT 1180.580000 0.000000 1181.980000 1.100000 ;
      RECT 1177.820000 0.000000 1179.680000 1.100000 ;
      RECT 1175.520000 0.000000 1176.920000 1.100000 ;
      RECT 1173.220000 0.000000 1174.620000 1.100000 ;
      RECT 1170.460000 0.000000 1172.320000 1.100000 ;
      RECT 1168.160000 0.000000 1169.560000 1.100000 ;
      RECT 1165.400000 0.000000 1167.260000 1.100000 ;
      RECT 1163.100000 0.000000 1164.500000 1.100000 ;
      RECT 1160.800000 0.000000 1162.200000 1.100000 ;
      RECT 1158.040000 0.000000 1159.900000 1.100000 ;
      RECT 1155.740000 0.000000 1157.140000 1.100000 ;
      RECT 1153.440000 0.000000 1154.840000 1.100000 ;
      RECT 1150.680000 0.000000 1152.540000 1.100000 ;
      RECT 1148.380000 0.000000 1149.780000 1.100000 ;
      RECT 1146.080000 0.000000 1147.480000 1.100000 ;
      RECT 1143.320000 0.000000 1145.180000 1.100000 ;
      RECT 1141.020000 0.000000 1142.420000 1.100000 ;
      RECT 1138.720000 0.000000 1140.120000 1.100000 ;
      RECT 1135.960000 0.000000 1137.820000 1.100000 ;
      RECT 1133.660000 0.000000 1135.060000 1.100000 ;
      RECT 1131.360000 0.000000 1132.760000 1.100000 ;
      RECT 1128.600000 0.000000 1130.460000 1.100000 ;
      RECT 1126.300000 0.000000 1127.700000 1.100000 ;
      RECT 1124.000000 0.000000 1125.400000 1.100000 ;
      RECT 1121.240000 0.000000 1123.100000 1.100000 ;
      RECT 1118.940000 0.000000 1120.340000 1.100000 ;
      RECT 1116.640000 0.000000 1118.040000 1.100000 ;
      RECT 1113.880000 0.000000 1115.740000 1.100000 ;
      RECT 1111.580000 0.000000 1112.980000 1.100000 ;
      RECT 1109.280000 0.000000 1110.680000 1.100000 ;
      RECT 1106.520000 0.000000 1108.380000 1.100000 ;
      RECT 1104.220000 0.000000 1105.620000 1.100000 ;
      RECT 1101.920000 0.000000 1103.320000 1.100000 ;
      RECT 1099.160000 0.000000 1101.020000 1.100000 ;
      RECT 1096.860000 0.000000 1098.260000 1.100000 ;
      RECT 1094.100000 0.000000 1095.960000 1.100000 ;
      RECT 1091.800000 0.000000 1093.200000 1.100000 ;
      RECT 1089.500000 0.000000 1090.900000 1.100000 ;
      RECT 1086.740000 0.000000 1088.600000 1.100000 ;
      RECT 1084.440000 0.000000 1085.840000 1.100000 ;
      RECT 1082.140000 0.000000 1083.540000 1.100000 ;
      RECT 1079.840000 0.000000 1081.240000 1.100000 ;
      RECT 1077.080000 0.000000 1078.940000 1.100000 ;
      RECT 1074.780000 0.000000 1076.180000 1.100000 ;
      RECT 1072.020000 0.000000 1073.880000 1.100000 ;
      RECT 1069.720000 0.000000 1071.120000 1.100000 ;
      RECT 1067.420000 0.000000 1068.820000 1.100000 ;
      RECT 1064.660000 0.000000 1066.520000 1.100000 ;
      RECT 1062.360000 0.000000 1063.760000 1.100000 ;
      RECT 1060.060000 0.000000 1061.460000 1.100000 ;
      RECT 1057.300000 0.000000 1059.160000 1.100000 ;
      RECT 1055.000000 0.000000 1056.400000 1.100000 ;
      RECT 1052.700000 0.000000 1054.100000 1.100000 ;
      RECT 1049.940000 0.000000 1051.800000 1.100000 ;
      RECT 1047.640000 0.000000 1049.040000 1.100000 ;
      RECT 1045.340000 0.000000 1046.740000 1.100000 ;
      RECT 1042.580000 0.000000 1044.440000 1.100000 ;
      RECT 1040.280000 0.000000 1041.680000 1.100000 ;
      RECT 1037.520000 0.000000 1039.380000 1.100000 ;
      RECT 1035.220000 0.000000 1036.620000 1.100000 ;
      RECT 1032.920000 0.000000 1034.320000 1.100000 ;
      RECT 1030.620000 0.000000 1032.020000 1.100000 ;
      RECT 1027.860000 0.000000 1029.720000 1.100000 ;
      RECT 1025.560000 0.000000 1026.960000 1.100000 ;
      RECT 1022.800000 0.000000 1024.660000 1.100000 ;
      RECT 1020.500000 0.000000 1021.900000 1.100000 ;
      RECT 1018.200000 0.000000 1019.600000 1.100000 ;
      RECT 1015.440000 0.000000 1017.300000 1.100000 ;
      RECT 1013.140000 0.000000 1014.540000 1.100000 ;
      RECT 1010.840000 0.000000 1012.240000 1.100000 ;
      RECT 1008.080000 0.000000 1009.940000 1.100000 ;
      RECT 1005.780000 0.000000 1007.180000 1.100000 ;
      RECT 1003.480000 0.000000 1004.880000 1.100000 ;
      RECT 1000.720000 0.000000 1002.580000 1.100000 ;
      RECT 998.420000 0.000000 999.820000 1.100000 ;
      RECT 996.120000 0.000000 997.520000 1.100000 ;
      RECT 993.360000 0.000000 995.220000 1.100000 ;
      RECT 991.060000 0.000000 992.460000 1.100000 ;
      RECT 988.300000 0.000000 990.160000 1.100000 ;
      RECT 986.000000 0.000000 987.400000 1.100000 ;
      RECT 983.700000 0.000000 985.100000 1.100000 ;
      RECT 981.400000 0.000000 982.800000 1.100000 ;
      RECT 978.640000 0.000000 980.500000 1.100000 ;
      RECT 976.340000 0.000000 977.740000 1.100000 ;
      RECT 974.040000 0.000000 975.440000 1.100000 ;
      RECT 971.280000 0.000000 973.140000 1.100000 ;
      RECT 968.980000 0.000000 970.380000 1.100000 ;
      RECT 966.680000 0.000000 968.080000 1.100000 ;
      RECT 963.920000 0.000000 965.780000 1.100000 ;
      RECT 961.620000 0.000000 963.020000 1.100000 ;
      RECT 959.320000 0.000000 960.720000 1.100000 ;
      RECT 956.560000 0.000000 958.420000 1.100000 ;
      RECT 954.260000 0.000000 955.660000 1.100000 ;
      RECT 951.500000 0.000000 953.360000 1.100000 ;
      RECT 949.200000 0.000000 950.600000 1.100000 ;
      RECT 946.900000 0.000000 948.300000 1.100000 ;
      RECT 944.140000 0.000000 946.000000 1.100000 ;
      RECT 941.840000 0.000000 943.240000 1.100000 ;
      RECT 939.540000 0.000000 940.940000 1.100000 ;
      RECT 936.780000 0.000000 938.640000 1.100000 ;
      RECT 934.480000 0.000000 935.880000 1.100000 ;
      RECT 932.180000 0.000000 933.580000 1.100000 ;
      RECT 929.420000 0.000000 931.280000 1.100000 ;
      RECT 927.120000 0.000000 928.520000 1.100000 ;
      RECT 924.820000 0.000000 926.220000 1.100000 ;
      RECT 922.060000 0.000000 923.920000 1.100000 ;
      RECT 919.760000 0.000000 921.160000 1.100000 ;
      RECT 917.460000 0.000000 918.860000 1.100000 ;
      RECT 914.700000 0.000000 916.560000 1.100000 ;
      RECT 912.400000 0.000000 913.800000 1.100000 ;
      RECT 910.100000 0.000000 911.500000 1.100000 ;
      RECT 907.340000 0.000000 909.200000 1.100000 ;
      RECT 905.040000 0.000000 906.440000 1.100000 ;
      RECT 902.740000 0.000000 904.140000 1.100000 ;
      RECT 899.980000 0.000000 901.840000 1.100000 ;
      RECT 897.680000 0.000000 899.080000 1.100000 ;
      RECT 894.920000 0.000000 896.780000 1.100000 ;
      RECT 892.620000 0.000000 894.020000 1.100000 ;
      RECT 890.320000 0.000000 891.720000 1.100000 ;
      RECT 887.560000 0.000000 889.420000 1.100000 ;
      RECT 885.260000 0.000000 886.660000 1.100000 ;
      RECT 882.960000 0.000000 884.360000 1.100000 ;
      RECT 880.200000 0.000000 882.060000 1.100000 ;
      RECT 877.900000 0.000000 879.300000 1.100000 ;
      RECT 875.600000 0.000000 877.000000 1.100000 ;
      RECT 872.840000 0.000000 874.700000 1.100000 ;
      RECT 870.540000 0.000000 871.940000 1.100000 ;
      RECT 868.240000 0.000000 869.640000 1.100000 ;
      RECT 865.480000 0.000000 867.340000 1.100000 ;
      RECT 863.180000 0.000000 864.580000 1.100000 ;
      RECT 860.880000 0.000000 862.280000 1.100000 ;
      RECT 858.120000 0.000000 859.980000 1.100000 ;
      RECT 855.820000 0.000000 857.220000 1.100000 ;
      RECT 853.520000 0.000000 854.920000 1.100000 ;
      RECT 850.760000 0.000000 852.620000 1.100000 ;
      RECT 848.460000 0.000000 849.860000 1.100000 ;
      RECT 846.160000 0.000000 847.560000 1.100000 ;
      RECT 843.400000 0.000000 845.260000 1.100000 ;
      RECT 841.100000 0.000000 842.500000 1.100000 ;
      RECT 838.800000 0.000000 840.200000 1.100000 ;
      RECT 836.040000 0.000000 837.900000 1.100000 ;
      RECT 833.740000 0.000000 835.140000 1.100000 ;
      RECT 831.440000 0.000000 832.840000 1.100000 ;
      RECT 828.680000 0.000000 830.540000 1.100000 ;
      RECT 826.380000 0.000000 827.780000 1.100000 ;
      RECT 823.620000 0.000000 825.480000 1.100000 ;
      RECT 821.320000 0.000000 822.720000 1.100000 ;
      RECT 819.020000 0.000000 820.420000 1.100000 ;
      RECT 816.720000 0.000000 818.120000 1.100000 ;
      RECT 813.960000 0.000000 815.820000 1.100000 ;
      RECT 811.660000 0.000000 813.060000 1.100000 ;
      RECT 808.900000 0.000000 810.760000 1.100000 ;
      RECT 806.600000 0.000000 808.000000 1.100000 ;
      RECT 804.300000 0.000000 805.700000 1.100000 ;
      RECT 801.540000 0.000000 803.400000 1.100000 ;
      RECT 799.240000 0.000000 800.640000 1.100000 ;
      RECT 796.940000 0.000000 798.340000 1.100000 ;
      RECT 794.180000 0.000000 796.040000 1.100000 ;
      RECT 791.880000 0.000000 793.280000 1.100000 ;
      RECT 789.580000 0.000000 790.980000 1.100000 ;
      RECT 786.820000 0.000000 788.680000 1.100000 ;
      RECT 784.520000 0.000000 785.920000 1.100000 ;
      RECT 782.220000 0.000000 783.620000 1.100000 ;
      RECT 779.460000 0.000000 781.320000 1.100000 ;
      RECT 777.160000 0.000000 778.560000 1.100000 ;
      RECT 774.400000 0.000000 776.260000 1.100000 ;
      RECT 772.100000 0.000000 773.500000 1.100000 ;
      RECT 769.800000 0.000000 771.200000 1.100000 ;
      RECT 767.500000 0.000000 768.900000 1.100000 ;
      RECT 764.740000 0.000000 766.600000 1.100000 ;
      RECT 762.440000 0.000000 763.840000 1.100000 ;
      RECT 760.140000 0.000000 761.540000 1.100000 ;
      RECT 757.380000 0.000000 759.240000 1.100000 ;
      RECT 755.080000 0.000000 756.480000 1.100000 ;
      RECT 752.320000 0.000000 754.180000 1.100000 ;
      RECT 750.020000 0.000000 751.420000 1.100000 ;
      RECT 747.720000 0.000000 749.120000 1.100000 ;
      RECT 744.960000 0.000000 746.820000 1.100000 ;
      RECT 742.660000 0.000000 744.060000 1.100000 ;
      RECT 740.360000 0.000000 741.760000 1.100000 ;
      RECT 737.600000 0.000000 739.460000 1.100000 ;
      RECT 735.300000 0.000000 736.700000 1.100000 ;
      RECT 733.000000 0.000000 734.400000 1.100000 ;
      RECT 730.240000 0.000000 732.100000 1.100000 ;
      RECT 727.940000 0.000000 729.340000 1.100000 ;
      RECT 725.640000 0.000000 727.040000 1.100000 ;
      RECT 722.880000 0.000000 724.740000 1.100000 ;
      RECT 720.580000 0.000000 721.980000 1.100000 ;
      RECT 718.280000 0.000000 719.680000 1.100000 ;
      RECT 715.520000 0.000000 717.380000 1.100000 ;
      RECT 713.220000 0.000000 714.620000 1.100000 ;
      RECT 710.920000 0.000000 712.320000 1.100000 ;
      RECT 708.160000 0.000000 710.020000 1.100000 ;
      RECT 705.860000 0.000000 707.260000 1.100000 ;
      RECT 703.560000 0.000000 704.960000 1.100000 ;
      RECT 700.800000 0.000000 702.660000 1.100000 ;
      RECT 698.500000 0.000000 699.900000 1.100000 ;
      RECT 696.200000 0.000000 697.600000 1.100000 ;
      RECT 693.440000 0.000000 695.300000 1.100000 ;
      RECT 691.140000 0.000000 692.540000 1.100000 ;
      RECT 688.840000 0.000000 690.240000 1.100000 ;
      RECT 686.080000 0.000000 687.940000 1.100000 ;
      RECT 683.780000 0.000000 685.180000 1.100000 ;
      RECT 681.020000 0.000000 682.880000 1.100000 ;
      RECT 678.720000 0.000000 680.120000 1.100000 ;
      RECT 676.420000 0.000000 677.820000 1.100000 ;
      RECT 673.660000 0.000000 675.520000 1.100000 ;
      RECT 671.360000 0.000000 672.760000 1.100000 ;
      RECT 669.060000 0.000000 670.460000 1.100000 ;
      RECT 666.300000 0.000000 668.160000 1.100000 ;
      RECT 664.000000 0.000000 665.400000 1.100000 ;
      RECT 661.700000 0.000000 663.100000 1.100000 ;
      RECT 658.940000 0.000000 660.800000 1.100000 ;
      RECT 656.640000 0.000000 658.040000 1.100000 ;
      RECT 654.340000 0.000000 655.740000 1.100000 ;
      RECT 651.580000 0.000000 653.440000 1.100000 ;
      RECT 649.280000 0.000000 650.680000 1.100000 ;
      RECT 646.980000 0.000000 648.380000 1.100000 ;
      RECT 644.220000 0.000000 646.080000 1.100000 ;
      RECT 641.920000 0.000000 643.320000 1.100000 ;
      RECT 639.620000 0.000000 641.020000 1.100000 ;
      RECT 636.860000 0.000000 638.720000 1.100000 ;
      RECT 634.560000 0.000000 635.960000 1.100000 ;
      RECT 631.800000 0.000000 633.660000 1.100000 ;
      RECT 629.500000 0.000000 630.900000 1.100000 ;
      RECT 627.200000 0.000000 628.600000 1.100000 ;
      RECT 624.440000 0.000000 626.300000 1.100000 ;
      RECT 622.140000 0.000000 623.540000 1.100000 ;
      RECT 619.840000 0.000000 621.240000 1.100000 ;
      RECT 617.540000 0.000000 618.940000 1.100000 ;
      RECT 614.780000 0.000000 616.640000 1.100000 ;
      RECT 612.480000 0.000000 613.880000 1.100000 ;
      RECT 609.720000 0.000000 611.580000 1.100000 ;
      RECT 607.420000 0.000000 608.820000 1.100000 ;
      RECT 605.120000 0.000000 606.520000 1.100000 ;
      RECT 602.820000 0.000000 604.220000 1.100000 ;
      RECT 600.060000 0.000000 601.920000 1.100000 ;
      RECT 597.760000 0.000000 599.160000 1.100000 ;
      RECT 595.000000 0.000000 596.860000 1.100000 ;
      RECT 592.700000 0.000000 594.100000 1.100000 ;
      RECT 590.400000 0.000000 591.800000 1.100000 ;
      RECT 587.640000 0.000000 589.500000 1.100000 ;
      RECT 585.340000 0.000000 586.740000 1.100000 ;
      RECT 583.040000 0.000000 584.440000 1.100000 ;
      RECT 580.280000 0.000000 582.140000 1.100000 ;
      RECT 577.980000 0.000000 579.380000 1.100000 ;
      RECT 575.680000 0.000000 577.080000 1.100000 ;
      RECT 572.920000 0.000000 574.780000 1.100000 ;
      RECT 570.620000 0.000000 572.020000 1.100000 ;
      RECT 568.320000 0.000000 569.720000 1.100000 ;
      RECT 565.560000 0.000000 567.420000 1.100000 ;
      RECT 563.260000 0.000000 564.660000 1.100000 ;
      RECT 560.500000 0.000000 562.360000 1.100000 ;
      RECT 558.200000 0.000000 559.600000 1.100000 ;
      RECT 555.900000 0.000000 557.300000 1.100000 ;
      RECT 553.600000 0.000000 555.000000 1.100000 ;
      RECT 550.840000 0.000000 552.700000 1.100000 ;
      RECT 548.540000 0.000000 549.940000 1.100000 ;
      RECT 546.240000 0.000000 547.640000 1.100000 ;
      RECT 543.480000 0.000000 545.340000 1.100000 ;
      RECT 541.180000 0.000000 542.580000 1.100000 ;
      RECT 538.420000 0.000000 540.280000 1.100000 ;
      RECT 536.120000 0.000000 537.520000 1.100000 ;
      RECT 533.820000 0.000000 535.220000 1.100000 ;
      RECT 531.060000 0.000000 532.920000 1.100000 ;
      RECT 528.760000 0.000000 530.160000 1.100000 ;
      RECT 526.460000 0.000000 527.860000 1.100000 ;
      RECT 523.700000 0.000000 525.560000 1.100000 ;
      RECT 521.400000 0.000000 522.800000 1.100000 ;
      RECT 519.100000 0.000000 520.500000 1.100000 ;
      RECT 516.340000 0.000000 518.200000 1.100000 ;
      RECT 514.040000 0.000000 515.440000 1.100000 ;
      RECT 511.740000 0.000000 513.140000 1.100000 ;
      RECT 508.980000 0.000000 510.840000 1.100000 ;
      RECT 506.680000 0.000000 508.080000 1.100000 ;
      RECT 504.380000 0.000000 505.780000 1.100000 ;
      RECT 501.620000 0.000000 503.480000 1.100000 ;
      RECT 499.320000 0.000000 500.720000 1.100000 ;
      RECT 497.020000 0.000000 498.420000 1.100000 ;
      RECT 494.260000 0.000000 496.120000 1.100000 ;
      RECT 491.960000 0.000000 493.360000 1.100000 ;
      RECT 489.660000 0.000000 491.060000 1.100000 ;
      RECT 486.900000 0.000000 488.760000 1.100000 ;
      RECT 484.600000 0.000000 486.000000 1.100000 ;
      RECT 482.300000 0.000000 483.700000 1.100000 ;
      RECT 479.540000 0.000000 481.400000 1.100000 ;
      RECT 477.240000 0.000000 478.640000 1.100000 ;
      RECT 474.940000 0.000000 476.340000 1.100000 ;
      RECT 472.180000 0.000000 474.040000 1.100000 ;
      RECT 469.880000 0.000000 471.280000 1.100000 ;
      RECT 467.120000 0.000000 468.980000 1.100000 ;
      RECT 464.820000 0.000000 466.220000 1.100000 ;
      RECT 462.520000 0.000000 463.920000 1.100000 ;
      RECT 459.760000 0.000000 461.620000 1.100000 ;
      RECT 457.460000 0.000000 458.860000 1.100000 ;
      RECT 455.160000 0.000000 456.560000 1.100000 ;
      RECT 452.400000 0.000000 454.260000 1.100000 ;
      RECT 450.100000 0.000000 451.500000 1.100000 ;
      RECT 447.800000 0.000000 449.200000 1.100000 ;
      RECT 445.040000 0.000000 446.900000 1.100000 ;
      RECT 442.740000 0.000000 444.140000 1.100000 ;
      RECT 440.440000 0.000000 441.840000 1.100000 ;
      RECT 437.680000 0.000000 439.540000 1.100000 ;
      RECT 435.380000 0.000000 436.780000 1.100000 ;
      RECT 433.080000 0.000000 434.480000 1.100000 ;
      RECT 430.320000 0.000000 432.180000 1.100000 ;
      RECT 428.020000 0.000000 429.420000 1.100000 ;
      RECT 425.720000 0.000000 427.120000 1.100000 ;
      RECT 422.960000 0.000000 424.820000 1.100000 ;
      RECT 420.660000 0.000000 422.060000 1.100000 ;
      RECT 417.900000 0.000000 419.760000 1.100000 ;
      RECT 415.600000 0.000000 417.000000 1.100000 ;
      RECT 413.300000 0.000000 414.700000 1.100000 ;
      RECT 410.540000 0.000000 412.400000 1.100000 ;
      RECT 408.240000 0.000000 409.640000 1.100000 ;
      RECT 405.940000 0.000000 407.340000 1.100000 ;
      RECT 403.640000 0.000000 405.040000 1.100000 ;
      RECT 400.880000 0.000000 402.740000 1.100000 ;
      RECT 398.580000 0.000000 399.980000 1.100000 ;
      RECT 395.820000 0.000000 397.680000 1.100000 ;
      RECT 393.520000 0.000000 394.920000 1.100000 ;
      RECT 391.220000 0.000000 392.620000 1.100000 ;
      RECT 388.460000 0.000000 390.320000 1.100000 ;
      RECT 386.160000 0.000000 387.560000 1.100000 ;
      RECT 383.860000 0.000000 385.260000 1.100000 ;
      RECT 381.100000 0.000000 382.960000 1.100000 ;
      RECT 378.800000 0.000000 380.200000 1.100000 ;
      RECT 376.500000 0.000000 377.900000 1.100000 ;
      RECT 373.740000 0.000000 375.600000 1.100000 ;
      RECT 371.440000 0.000000 372.840000 1.100000 ;
      RECT 369.140000 0.000000 370.540000 1.100000 ;
      RECT 366.380000 0.000000 368.240000 1.100000 ;
      RECT 364.080000 0.000000 365.480000 1.100000 ;
      RECT 361.780000 0.000000 363.180000 1.100000 ;
      RECT 359.020000 0.000000 360.880000 1.100000 ;
      RECT 356.720000 0.000000 358.120000 1.100000 ;
      RECT 354.420000 0.000000 355.820000 1.100000 ;
      RECT 351.660000 0.000000 353.520000 1.100000 ;
      RECT 349.360000 0.000000 350.760000 1.100000 ;
      RECT 346.600000 0.000000 348.460000 1.100000 ;
      RECT 344.300000 0.000000 345.700000 1.100000 ;
      RECT 342.000000 0.000000 343.400000 1.100000 ;
      RECT 339.700000 0.000000 341.100000 1.100000 ;
      RECT 336.940000 0.000000 338.800000 1.100000 ;
      RECT 334.640000 0.000000 336.040000 1.100000 ;
      RECT 332.340000 0.000000 333.740000 1.100000 ;
      RECT 329.580000 0.000000 331.440000 1.100000 ;
      RECT 327.280000 0.000000 328.680000 1.100000 ;
      RECT 324.520000 0.000000 326.380000 1.100000 ;
      RECT 322.220000 0.000000 323.620000 1.100000 ;
      RECT 319.920000 0.000000 321.320000 1.100000 ;
      RECT 317.160000 0.000000 319.020000 1.100000 ;
      RECT 314.860000 0.000000 316.260000 1.100000 ;
      RECT 312.560000 0.000000 313.960000 1.100000 ;
      RECT 309.800000 0.000000 311.660000 1.100000 ;
      RECT 307.500000 0.000000 308.900000 1.100000 ;
      RECT 305.200000 0.000000 306.600000 1.100000 ;
      RECT 302.440000 0.000000 304.300000 1.100000 ;
      RECT 300.140000 0.000000 301.540000 1.100000 ;
      RECT 297.840000 0.000000 299.240000 1.100000 ;
      RECT 295.080000 0.000000 296.940000 1.100000 ;
      RECT 292.780000 0.000000 294.180000 1.100000 ;
      RECT 290.480000 0.000000 291.880000 1.100000 ;
      RECT 287.720000 0.000000 289.580000 1.100000 ;
      RECT 285.420000 0.000000 286.820000 1.100000 ;
      RECT 283.120000 0.000000 284.520000 1.100000 ;
      RECT 280.360000 0.000000 282.220000 1.100000 ;
      RECT 278.060000 0.000000 279.460000 1.100000 ;
      RECT 275.300000 0.000000 277.160000 1.100000 ;
      RECT 273.000000 0.000000 274.400000 1.100000 ;
      RECT 270.700000 0.000000 272.100000 1.100000 ;
      RECT 267.940000 0.000000 269.800000 1.100000 ;
      RECT 265.640000 0.000000 267.040000 1.100000 ;
      RECT 263.340000 0.000000 264.740000 1.100000 ;
      RECT 260.580000 0.000000 262.440000 1.100000 ;
      RECT 258.280000 0.000000 259.680000 1.100000 ;
      RECT 255.980000 0.000000 257.380000 1.100000 ;
      RECT 253.220000 0.000000 255.080000 1.100000 ;
      RECT 250.920000 0.000000 252.320000 1.100000 ;
      RECT 248.620000 0.000000 250.020000 1.100000 ;
      RECT 245.860000 0.000000 247.720000 1.100000 ;
      RECT 243.560000 0.000000 244.960000 1.100000 ;
      RECT 241.260000 0.000000 242.660000 1.100000 ;
      RECT 238.500000 0.000000 240.360000 1.100000 ;
      RECT 236.200000 0.000000 237.600000 1.100000 ;
      RECT 233.900000 0.000000 235.300000 1.100000 ;
      RECT 231.140000 0.000000 233.000000 1.100000 ;
      RECT 228.840000 0.000000 230.240000 1.100000 ;
      RECT 226.540000 0.000000 227.940000 1.100000 ;
      RECT 223.780000 0.000000 225.640000 1.100000 ;
      RECT 221.480000 0.000000 222.880000 1.100000 ;
      RECT 219.180000 0.000000 220.580000 1.100000 ;
      RECT 216.420000 0.000000 218.280000 1.100000 ;
      RECT 214.120000 0.000000 215.520000 1.100000 ;
      RECT 211.820000 0.000000 213.220000 1.100000 ;
      RECT 209.060000 0.000000 210.920000 1.100000 ;
      RECT 206.760000 0.000000 208.160000 1.100000 ;
      RECT 204.000000 0.000000 205.860000 1.100000 ;
      RECT 201.700000 0.000000 203.100000 1.100000 ;
      RECT 199.400000 0.000000 200.800000 1.100000 ;
      RECT 196.640000 0.000000 198.500000 1.100000 ;
      RECT 194.340000 0.000000 195.740000 1.100000 ;
      RECT 192.040000 0.000000 193.440000 1.100000 ;
      RECT 189.740000 0.000000 191.140000 1.100000 ;
      RECT 186.980000 0.000000 188.840000 1.100000 ;
      RECT 184.680000 0.000000 186.080000 1.100000 ;
      RECT 181.920000 0.000000 183.780000 1.100000 ;
      RECT 179.620000 0.000000 181.020000 1.100000 ;
      RECT 177.320000 0.000000 178.720000 1.100000 ;
      RECT 174.560000 0.000000 176.420000 1.100000 ;
      RECT 172.260000 0.000000 173.660000 1.100000 ;
      RECT 169.960000 0.000000 171.360000 1.100000 ;
      RECT 167.200000 0.000000 169.060000 1.100000 ;
      RECT 164.900000 0.000000 166.300000 1.100000 ;
      RECT 162.600000 0.000000 164.000000 1.100000 ;
      RECT 159.840000 0.000000 161.700000 1.100000 ;
      RECT 157.540000 0.000000 158.940000 1.100000 ;
      RECT 155.240000 0.000000 156.640000 1.100000 ;
      RECT 152.480000 0.000000 154.340000 1.100000 ;
      RECT 150.180000 0.000000 151.580000 1.100000 ;
      RECT 147.420000 0.000000 149.280000 1.100000 ;
      RECT 145.120000 0.000000 146.520000 1.100000 ;
      RECT 142.820000 0.000000 144.220000 1.100000 ;
      RECT 140.520000 0.000000 141.920000 1.100000 ;
      RECT 137.760000 0.000000 139.620000 1.100000 ;
      RECT 135.460000 0.000000 136.860000 1.100000 ;
      RECT 132.700000 0.000000 134.560000 1.100000 ;
      RECT 130.400000 0.000000 131.800000 1.100000 ;
      RECT 128.100000 0.000000 129.500000 1.100000 ;
      RECT 125.800000 0.000000 127.200000 1.100000 ;
      RECT 123.040000 0.000000 124.900000 1.100000 ;
      RECT 120.740000 0.000000 122.140000 1.100000 ;
      RECT 118.440000 0.000000 119.840000 1.100000 ;
      RECT 115.680000 0.000000 117.540000 1.100000 ;
      RECT 113.380000 0.000000 114.780000 1.100000 ;
      RECT 110.620000 0.000000 112.480000 1.100000 ;
      RECT 108.320000 0.000000 109.720000 1.100000 ;
      RECT 106.020000 0.000000 107.420000 1.100000 ;
      RECT 103.260000 0.000000 105.120000 1.100000 ;
      RECT 100.960000 0.000000 102.360000 1.100000 ;
      RECT 98.660000 0.000000 100.060000 1.100000 ;
      RECT 95.900000 0.000000 97.760000 1.100000 ;
      RECT 93.600000 0.000000 95.000000 1.100000 ;
      RECT 91.300000 0.000000 92.700000 1.100000 ;
      RECT 88.540000 0.000000 90.400000 1.100000 ;
      RECT 86.240000 0.000000 87.640000 1.100000 ;
      RECT 83.940000 0.000000 85.340000 1.100000 ;
      RECT 81.180000 0.000000 83.040000 1.100000 ;
      RECT 78.880000 0.000000 80.280000 1.100000 ;
      RECT 76.580000 0.000000 77.980000 1.100000 ;
      RECT 73.820000 0.000000 75.680000 1.100000 ;
      RECT 71.520000 0.000000 72.920000 1.100000 ;
      RECT 69.220000 0.000000 70.620000 1.100000 ;
      RECT 66.460000 0.000000 68.320000 1.100000 ;
      RECT 64.160000 0.000000 65.560000 1.100000 ;
      RECT 61.400000 0.000000 63.260000 1.100000 ;
      RECT 59.100000 0.000000 60.500000 1.100000 ;
      RECT 56.800000 0.000000 58.200000 1.100000 ;
      RECT 54.040000 0.000000 55.900000 1.100000 ;
      RECT 51.740000 0.000000 53.140000 1.100000 ;
      RECT 49.440000 0.000000 50.840000 1.100000 ;
      RECT 46.680000 0.000000 48.540000 1.100000 ;
      RECT 44.380000 0.000000 45.780000 1.100000 ;
      RECT 42.080000 0.000000 43.480000 1.100000 ;
      RECT 39.320000 0.000000 41.180000 1.100000 ;
      RECT 37.020000 0.000000 38.420000 1.100000 ;
      RECT 34.720000 0.000000 36.120000 1.100000 ;
      RECT 31.960000 0.000000 33.820000 1.100000 ;
      RECT 29.660000 0.000000 31.060000 1.100000 ;
      RECT 27.360000 0.000000 28.760000 1.100000 ;
      RECT 24.600000 0.000000 26.460000 1.100000 ;
      RECT 22.300000 0.000000 23.700000 1.100000 ;
      RECT 20.000000 0.000000 21.400000 1.100000 ;
      RECT 17.240000 0.000000 19.100000 1.100000 ;
      RECT 14.940000 0.000000 16.340000 1.100000 ;
      RECT 12.640000 0.000000 14.040000 1.100000 ;
      RECT 9.880000 0.000000 11.740000 1.100000 ;
      RECT 7.580000 0.000000 8.980000 1.100000 ;
      RECT 4.820000 0.000000 6.680000 1.100000 ;
      RECT 2.520000 0.000000 3.920000 1.100000 ;
      RECT 1.600000 0.000000 1.620000 1.100000 ;
      RECT 0.000000 0.000000 0.700000 0.180000 ;
    LAYER met4 ;
      RECT 0.000000 1056.620000 1222.220000 1061.140000 ;
      RECT 6.540000 1053.420000 1215.680000 1056.620000 ;
      RECT 1214.680000 7.380000 1215.680000 1053.420000 ;
      RECT 9.740000 7.380000 1212.480000 1053.420000 ;
      RECT 6.540000 7.380000 7.540000 1053.420000 ;
      RECT 1217.880000 4.180000 1222.220000 1056.620000 ;
      RECT 6.540000 4.180000 1215.680000 7.380000 ;
      RECT 0.000000 4.180000 4.340000 1056.620000 ;
      RECT 0.000000 0.000000 1222.220000 4.180000 ;
  END
END soc_now_caravel_top

END LIBRARY
